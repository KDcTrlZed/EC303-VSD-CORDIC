* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : cordic_pipeline                              *
* Netlisted  : Mon Oct 21 14:42:59 2024                     *
* PVS Version: 22.20-p031 Thu Nov 17 19:06:38 PST 2022      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(nmos1v) _nmos_12 ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(pmos1v) _pmos_12 pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: CLKBUFX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt CLKBUFX2 Y VDD VSS A
** N=5 EP=4 FDC=6
M0 Y 5 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=830 $dt=0
M1 VSS 5 Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1550 $Y=830 $dt=0
M2 5 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2390 $Y=1060 $dt=0
M3 Y 5 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=2940 $dt=1
M4 VDD 5 Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1550 $Y=2940 $dt=1
M5 5 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2390 $Y=3000 $dt=1
.ends CLKBUFX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: CLKINVX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt CLKINVX2 A VDD VSS Y
** N=4 EP=4 FDC=4
M0 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=900 $Y=980 $dt=0
M1 VSS A Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1740 $Y=980 $dt=0
M2 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=900 $Y=2720 $dt=1
M3 VDD A Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1740 $Y=2720 $dt=1
.ends CLKINVX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: CLKINVX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt CLKINVX1 A Y VDD VSS
** N=4 EP=4 FDC=2
M0 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=870 $dt=0
M1 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=2680 $dt=1
.ends CLKINVX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFFRHQX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFFRHQX1 Q CK VDD VSS RN D
** N=20 EP=6 FDC=28
M0 VSS 11 Q VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=900 $dt=0
M1 7 CK VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1790 $Y=1230 $dt=0
M2 13 12 11 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=3430 $Y=800 $dt=0
M3 VSS RN 13 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=3870 $Y=800 $dt=0
M4 14 11 VSS VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=5150 $Y=800 $dt=0
M5 12 7 14 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=5870 $Y=800 $dt=0
M6 9 8 12 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=7390 $Y=880 $dt=0
M7 VSS 10 9 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=8350 $Y=880 $dt=0
M8 15 RN VSS VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=9670 $Y=880 $dt=0
M9 16 9 15 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=10110 $Y=880 $dt=0
M10 10 8 16 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=11030 $Y=880 $dt=0
M11 17 7 10 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=11870 $Y=880 $dt=0
M12 VSS D 17 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=12310 $Y=880 $dt=0
M13 8 7 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=14630 $Y=800 $dt=0
M14 VDD 11 Q VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=2680 $dt=1
M15 7 CK VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=3000 $dt=1
M16 11 12 VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=3430 $Y=3080 $dt=1
M17 VDD RN 11 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=4270 $Y=3080 $dt=1
M18 19 11 VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=5510 $Y=2940 $dt=1
M19 12 8 19 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=5950 $Y=2940 $dt=1
M20 9 7 12 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=6910 $Y=2940 $dt=1
M21 VDD 10 9 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=7750 $Y=2940 $dt=1
M22 18 RN VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=9150 $Y=2940 $dt=1
M23 VDD 9 18 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=9990 $Y=3380 $dt=1
M24 10 7 18 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=11990 $Y=3040 $dt=1
M25 20 8 10 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=12950 $Y=3340 $dt=1
M26 VDD D 20 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=13550 $Y=3340 $dt=1
M27 8 7 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=14630 $Y=3140 $dt=1
.ends DFFRHQX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: SDFFRHQX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt SDFFRHQX1 Q CK VDD VSS RN D SI SE
** N=26 EP=8 FDC=36
M0 VSS 14 Q VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=980 $dt=0
M1 10 CK VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1670 $Y=1360 $dt=0
M2 16 15 14 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=3410 $Y=880 $dt=0
M3 VSS RN 16 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=4170 $Y=880 $dt=0
M4 17 14 VSS VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=5250 $Y=880 $dt=0
M5 15 10 17 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=5890 $Y=880 $dt=0
M6 12 11 15 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=7570 $Y=880 $dt=0
M7 VSS 13 12 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=8690 $Y=880 $dt=0
M8 18 RN VSS VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=9930 $Y=880 $dt=0
M9 19 12 18 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=10370 $Y=880 $dt=0
M10 13 11 19 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=10810 $Y=880 $dt=0
M11 20 10 13 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=11650 $Y=880 $dt=0
M12 VSS 10 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=14090 $Y=1180 $dt=0
M13 21 D VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=15050 $Y=800 $dt=0
M14 20 9 21 VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=16010 $Y=800 $dt=0
M15 22 SE 20 VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=16850 $Y=800 $dt=0
M16 VSS SI 22 VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=17290 $Y=800 $dt=0
M17 9 SE VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=18130 $Y=1160 $dt=0
M18 VDD 14 Q VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=2720 $dt=1
M19 10 CK VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=3110 $dt=1
M20 14 15 VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=3410 $Y=2940 $dt=1
M21 VDD RN 14 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=4330 $Y=2940 $dt=1
M22 23 14 VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=5450 $Y=2940 $dt=1
M23 15 11 23 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=5890 $Y=2940 $dt=1
M24 12 10 15 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=6850 $Y=2940 $dt=1
M25 VDD 13 12 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=7810 $Y=2940 $dt=1
M26 24 RN VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=9130 $Y=2940 $dt=1
M27 VDD 12 24 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=9970 $Y=2940 $dt=1
M28 13 10 24 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=11710 $Y=2840 $dt=1
M29 20 11 13 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=12550 $Y=2840 $dt=1
M30 VDD 10 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=14170 $Y=3120 $dt=1
M31 25 D VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=15050 $Y=3120 $dt=1
M32 20 SE 25 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=15490 $Y=3120 $dt=1
M33 26 9 20 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=16330 $Y=3120 $dt=1
M34 VDD SI 26 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=16970 $Y=3120 $dt=1
M35 9 SE VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=18010 $Y=3120 $dt=1
.ends SDFFRHQX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFFRX1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFFRX1 QN VDD VSS Q CK RN D
** N=22 EP=7 FDC=32
M0 VSS 14 QN VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=980 $dt=0
M1 14 12 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1570 $Y=1360 $dt=0
M2 VSS 12 Q VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=3190 $Y=840 $dt=0
M3 8 CK VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4270 $Y=1220 $dt=0
M4 15 13 12 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5910 $Y=1100 $dt=0
M5 VSS RN 15 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=6350 $Y=1100 $dt=0
M6 16 12 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7730 $Y=1100 $dt=0
M7 13 8 16 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=8170 $Y=1100 $dt=0
M8 10 9 13 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=9070 $Y=1100 $dt=0
M9 VSS 11 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=10210 $Y=1100 $dt=0
M10 17 RN VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=11530 $Y=1240 $dt=0
M11 18 10 17 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=12030 $Y=1240 $dt=0
M12 11 9 18 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=12690 $Y=1240 $dt=0
M13 19 8 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=13530 $Y=1240 $dt=0
M14 VSS D 19 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=13970 $Y=1240 $dt=0
M15 9 8 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=15250 $Y=1240 $dt=0
M16 VDD 14 QN VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=2680 $dt=1
M17 14 12 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=2680 $dt=1
M18 VDD 12 Q VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=3010 $Y=3120 $dt=1
M19 8 CK VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3850 $Y=3120 $dt=1
M20 12 13 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5510 $Y=3020 $dt=1
M21 VDD RN 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=6350 $Y=3020 $dt=1
M22 20 12 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7350 $Y=3020 $dt=1
M23 13 9 20 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7790 $Y=3020 $dt=1
M24 10 8 13 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=8630 $Y=3020 $dt=1
M25 VDD 11 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=10230 $Y=3020 $dt=1
M26 21 RN VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=11190 $Y=3020 $dt=1
M27 VDD 10 21 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=12030 $Y=3020 $dt=1
M28 11 8 21 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=13530 $Y=3260 $dt=1
M29 22 9 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=14370 $Y=3260 $dt=1
M30 VDD D 22 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=14810 $Y=3260 $dt=1
M31 9 8 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=15890 $Y=3140 $dt=1
.ends DFFRX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: SDFFRXL                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt SDFFRXL QN VDD VSS Q CK RN D SE SI
** N=28 EP=9 FDC=40
M0 VSS 17 QN VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1360 $dt=0
M1 17 15 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1570 $Y=1360 $dt=0
M2 VSS 15 Q VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3190 $Y=1360 $dt=0
M3 11 CK VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4110 $Y=1360 $dt=0
M4 18 16 15 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5750 $Y=1240 $dt=0
M5 VSS RN 18 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=6190 $Y=1240 $dt=0
M6 19 15 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7270 $Y=1240 $dt=0
M7 16 11 19 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7910 $Y=1240 $dt=0
M8 13 12 16 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=9230 $Y=1240 $dt=0
M9 VSS 14 13 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=10310 $Y=1240 $dt=0
M10 20 RN VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=11390 $Y=1240 $dt=0
M11 21 13 20 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=11830 $Y=1240 $dt=0
M12 14 12 21 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=12550 $Y=1240 $dt=0
M13 22 11 14 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=13390 $Y=1240 $dt=0
M14 VSS 11 12 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=15550 $Y=800 $dt=0
M15 23 D VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=16510 $Y=800 $dt=0
M16 22 10 23 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=17390 $Y=800 $dt=0
M17 24 SE 22 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=18230 $Y=800 $dt=0
M18 VSS SI 24 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=18670 $Y=800 $dt=0
M19 10 SE VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=19510 $Y=800 $dt=0
M20 VDD 17 QN VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=2680 $dt=1
M21 17 15 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1790 $Y=2680 $dt=1
M22 VDD 15 Q VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3110 $Y=3700 $dt=1
M23 11 CK VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3950 $Y=3700 $dt=1
M24 15 16 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5690 $Y=3020 $dt=1
M25 VDD RN 15 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=6530 $Y=3020 $dt=1
M26 25 15 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7550 $Y=3020 $dt=1
M27 16 12 25 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7990 $Y=3020 $dt=1
M28 13 11 16 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=9150 $Y=3020 $dt=1
M29 VDD 14 13 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=10030 $Y=3020 $dt=1
M30 26 RN VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=10870 $Y=3020 $dt=1
M31 VDD 13 26 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=11710 $Y=3020 $dt=1
M32 14 11 26 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=13210 $Y=2720 $dt=1
M33 22 12 14 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=14050 $Y=2720 $dt=1
M34 VDD 11 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=15670 $Y=2880 $dt=1
M35 27 D VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=16510 $Y=2880 $dt=1
M36 22 SE 27 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=16950 $Y=2880 $dt=1
M37 28 10 22 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=17790 $Y=2880 $dt=1
M38 VDD SI 28 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=18670 $Y=2880 $dt=1
M39 10 SE VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=19510 $Y=2880 $dt=1
.ends SDFFRXL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XNOR3X1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XNOR3X1 A B VDD VSS C Y
** N=13 EP=6 FDC=22
M0 VSS A 11 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=970 $Y=800 $dt=0
M1 10 B VSS VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=2050 $Y=800 $dt=0
M2 9 11 VSS VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=4410 $Y=800 $dt=0
M3 12 B 9 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=5490 $Y=800 $dt=0
M4 11 10 12 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=7270 $Y=800 $dt=0
M5 13 B 11 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=8680 $Y=800 $dt=0
M6 9 10 13 VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=9760 $Y=800 $dt=0
M7 7 C 12 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=12120 $Y=800 $dt=0
M8 13 8 7 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=13200 $Y=800 $dt=0
M9 VSS C 8 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=15060 $Y=800 $dt=0
M10 Y 7 VSS VSS nmos1v L=1e-07 W=3.4e-07 fw=3.4e-07 simw=3.4e-07 $X=16140 $Y=800 $dt=0
M11 VDD A 11 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=970 $Y=3120 $dt=1
M12 10 B VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=2050 $Y=3380 $dt=1
M13 9 11 VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=4410 $Y=3380 $dt=1
M14 12 10 9 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=5490 $Y=3380 $dt=1
M15 11 B 12 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=6650 $Y=3080 $dt=1
M16 13 10 11 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=8150 $Y=2680 $dt=1
M17 9 B 13 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=9750 $Y=3340 $dt=1
M18 7 8 12 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=12120 $Y=3380 $dt=1
M19 13 C 7 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=13200 $Y=3380 $dt=1
M20 VDD C 8 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=15060 $Y=3380 $dt=1
M21 Y 7 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=16140 $Y=3120 $dt=1
.ends XNOR3X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OAI221XL                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OAI221XL A0 VDD VSS A1 B1 Y B0 C0
** N=12 EP=8 FDC=10
M0 9 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=640 $Y=1320 $dt=0
M1 VSS A1 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1480 $Y=1320 $dt=0
M2 9 B1 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2980 $Y=1360 $dt=0
M3 10 B0 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3820 $Y=1360 $dt=0
M4 Y C0 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4660 $Y=1360 $dt=0
M5 11 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1040 $Y=3410 $dt=1
M6 Y A1 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1480 $Y=3410 $dt=1
M7 12 B1 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2480 $Y=3410 $dt=1
M8 VDD B0 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2920 $Y=3410 $dt=1
M9 Y C0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4180 $Y=3410 $dt=1
.ends OAI221XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR3X1                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR3X1 C B VDD VSS A Y
** N=9 EP=6 FDC=8
M0 VSS C 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=800 $dt=0
M1 7 B VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1550 $Y=800 $dt=0
M2 VSS A 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2390 $Y=800 $dt=0
M3 Y 7 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=3230 $Y=800 $dt=0
M4 8 C 7 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=870 $Y=2850 $dt=1
M5 9 B 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=2850 $dt=1
M6 VDD A 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2230 $Y=2850 $dt=1
M7 Y 7 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=3190 $Y=2680 $dt=1
.ends OR3X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OAI211XL                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OAI211XL A0 VDD VSS Y A1 B0 C0
** N=10 EP=7 FDC=8
M0 VSS A0 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1140 $dt=0
M1 8 A1 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1550 $Y=1140 $dt=0
M2 9 B0 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2390 $Y=1140 $dt=0
M3 Y C0 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2830 $Y=1140 $dt=0
M4 10 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=820 $Y=3180 $dt=1
M5 Y A1 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1260 $Y=3180 $dt=1
M6 VDD B0 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2100 $Y=3180 $dt=1
M7 Y C0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3150 $Y=3180 $dt=1
.ends OAI211XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OAI32XL                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OAI32XL A0 VDD VSS A1 A2 Y B1 B0
** N=12 EP=8 FDC=10
M0 9 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=840 $Y=1270 $dt=0
M1 VSS A1 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1680 $Y=1270 $dt=0
M2 9 A2 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2520 $Y=1270 $dt=0
M3 Y B1 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3360 $Y=1270 $dt=0
M4 9 B0 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4200 $Y=1270 $dt=0
M5 10 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=840 $Y=3510 $dt=1
M6 11 A1 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1680 $Y=3510 $dt=1
M7 Y A2 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2520 $Y=3510 $dt=1
M8 12 B1 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3610 $Y=3510 $dt=1
M9 VDD B0 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4250 $Y=3510 $dt=1
.ends OAI32XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR2X1                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR2X1 B VDD VSS A Y
** N=7 EP=5 FDC=6
M0 6 B VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=770 $Y=1320 $dt=0
M1 VSS A 6 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1610 $Y=1320 $dt=0
M2 Y 6 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=2570 $Y=940 $dt=0
M3 7 B 6 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1170 $Y=3100 $dt=1
M4 VDD A 7 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1610 $Y=3100 $dt=1
M5 Y 6 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=2570 $Y=3100 $dt=1
.ends OR2X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NOR2BXL                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NOR2BXL Y B VDD VSS AN
** N=7 EP=5 FDC=6
M0 Y B VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=800 $dt=0
M1 VSS 6 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1550 $Y=800 $dt=0
M2 6 AN VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2390 $Y=800 $dt=0
M3 7 B Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1110 $Y=2980 $dt=1
M4 VDD 6 7 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=2980 $dt=1
M5 6 AN VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2390 $Y=2980 $dt=1
.ends NOR2BXL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OA21X1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OA21X1 A0 A1 VDD VSS B0 Y
** N=9 EP=6 FDC=8
M0 VSS A0 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1360 $dt=0
M1 8 A1 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1580 $Y=1360 $dt=0
M2 7 B0 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2580 $Y=1360 $dt=0
M3 Y 7 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=4100 $Y=800 $dt=0
M4 9 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1140 $Y=3120 $dt=1
M5 7 A1 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1580 $Y=3120 $dt=1
M6 VDD B0 7 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2580 $Y=3120 $dt=1
M7 Y 7 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=3540 $Y=3120 $dt=1
.ends OA21X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MXI2XL                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MXI2XL A Y VDD VSS S0 B
** N=11 EP=6 FDC=10
M0 8 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=720 $Y=1320 $dt=0
M1 Y 7 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1160 $Y=1320 $dt=0
M2 9 S0 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2000 $Y=1320 $dt=0
M3 VSS B 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2460 $Y=1320 $dt=0
M4 7 S0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3300 $Y=1320 $dt=0
M5 10 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=720 $Y=3700 $dt=1
M6 Y S0 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1160 $Y=3700 $dt=1
M7 11 7 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2000 $Y=3700 $dt=1
M8 VDD B 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2440 $Y=3700 $dt=1
M9 7 S0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3280 $Y=3700 $dt=1
.ends MXI2XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND3X1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND3X1 C B VDD VSS A Y
** N=9 EP=6 FDC=8
M0 8 C 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=980 $Y=1360 $dt=0
M1 9 B 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1780 $Y=1360 $dt=0
M2 VSS A 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2260 $Y=1360 $dt=0
M3 Y 7 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=3220 $Y=980 $dt=0
M4 VDD C 7 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=3150 $dt=1
M5 7 B VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1780 $Y=3150 $dt=1
M6 VDD A 7 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2620 $Y=3150 $dt=1
M7 Y 7 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=3460 $Y=2720 $dt=1
.ends AND3X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AOI221XL                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AOI221XL A0 VDD VSS A1 B1 Y B0 C0
** N=12 EP=8 FDC=10
M0 9 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1070 $Y=800 $dt=0
M1 Y A1 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1510 $Y=800 $dt=0
M2 10 B1 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3050 $Y=800 $dt=0
M3 VSS B0 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3490 $Y=800 $dt=0
M4 Y C0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4330 $Y=800 $dt=0
M5 12 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=670 $Y=3180 $dt=1
M6 VDD A1 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1510 $Y=3180 $dt=1
M7 12 B1 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3050 $Y=2840 $dt=1
M8 11 B0 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3890 $Y=2840 $dt=1
M9 Y C0 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4730 $Y=2840 $dt=1
.ends AOI221XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BMXIX2                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BMXIX2 M0 S VDD VSS A M1 X2 PPN
** N=22 EP=8 FDC=30
M0 VSS M0 12 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1220 $dt=0
M1 13 S VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1550 $Y=1220 $dt=0
M2 14 12 13 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1990 $Y=1220 $dt=0
M3 15 M0 14 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2830 $Y=1220 $dt=0
M4 VSS A 15 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3270 $Y=1220 $dt=0
M5 16 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4990 $Y=1220 $dt=0
M6 17 M1 16 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5430 $Y=1220 $dt=0
M7 18 11 17 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=6270 $Y=1220 $dt=0
M8 VSS S 18 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=6710 $Y=1220 $dt=0
M9 11 M1 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7790 $Y=1240 $dt=0
M10 9 X2 14 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=9630 $Y=1260 $dt=0
M11 17 10 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=10470 $Y=1260 $dt=0
M12 VSS X2 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=12090 $Y=1340 $dt=0
M13 PPN 9 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=13170 $Y=960 $dt=0
M14 VSS 9 PPN VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=14010 $Y=960 $dt=0
M15 VDD M0 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1030 $Y=3460 $dt=1
M16 19 S VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1870 $Y=3460 $dt=1
M17 14 M0 19 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2310 $Y=3460 $dt=1
M18 20 12 14 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3150 $Y=3460 $dt=1
M19 VDD A 20 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3590 $Y=3460 $dt=1
M20 21 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4670 $Y=3460 $dt=1
M21 17 11 21 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5110 $Y=3460 $dt=1
M22 22 M1 17 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5950 $Y=3220 $dt=1
M23 VDD S 22 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=6710 $Y=3220 $dt=1
M24 11 M1 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7790 $Y=3020 $dt=1
M25 9 10 14 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=9590 $Y=3060 $dt=1
M26 17 X2 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=10470 $Y=3060 $dt=1
M27 VDD X2 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=12320 $Y=3060 $dt=1
M28 PPN 9 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=13160 $Y=2680 $dt=1
M29 VDD 9 PPN VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=14000 $Y=2680 $dt=1
.ends BMXIX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ADDHX1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ADDHX1 CO A VDD VSS B S
** N=13 EP=6 FDC=18
M0 VSS 10 CO VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=780 $Y=820 $dt=0
M1 11 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1740 $Y=1200 $dt=0
M2 10 B 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2180 $Y=1200 $dt=0
M3 VSS B 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4040 $Y=1240 $dt=0
M4 8 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5120 $Y=1240 $dt=0
M5 7 9 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5960 $Y=1240 $dt=0
M6 12 B 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=6800 $Y=1240 $dt=0
M7 VSS 8 12 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7480 $Y=1240 $dt=0
M8 S 7 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=8320 $Y=980 $dt=0
M9 VDD 10 CO VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=780 $Y=3120 $dt=1
M10 10 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1620 $Y=3700 $dt=1
M11 VDD B 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2460 $Y=3700 $dt=1
M12 VDD B 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4040 $Y=3260 $dt=1
M13 8 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5120 $Y=3260 $dt=1
M14 7 B 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=6200 $Y=3260 $dt=1
M15 13 9 7 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7040 $Y=3260 $dt=1
M16 VDD 8 13 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7480 $Y=3260 $dt=1
M17 S 7 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=8320 $Y=2680 $dt=1
.ends ADDHX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO21X1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO21X1 A0 VDD VSS A1 B0 Y
** N=9 EP=6 FDC=8
M0 8 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=960 $Y=800 $dt=0
M1 7 A1 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1600 $Y=800 $dt=0
M2 VSS B0 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2440 $Y=800 $dt=0
M3 Y 7 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=3280 $Y=800 $dt=0
M4 VDD A0 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=760 $Y=3000 $dt=1
M5 9 A1 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1600 $Y=3000 $dt=1
M6 7 B0 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2440 $Y=3000 $dt=1
M7 Y 7 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=3900 $Y=3120 $dt=1
.ends AO21X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XNOR2X1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XNOR2X1 Y A VDD VSS B
** N=10 EP=5 FDC=12
M0 VSS 8 Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1110 $Y=980 $dt=0
M1 6 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1950 $Y=1240 $dt=0
M2 8 B 6 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2790 $Y=1240 $dt=0
M3 9 7 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3630 $Y=1240 $dt=0
M4 VSS 6 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4630 $Y=1240 $dt=0
M5 7 B VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5470 $Y=1240 $dt=0
M6 VDD 8 Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=3080 $dt=1
M7 6 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=3080 $dt=1
M8 8 7 6 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2390 $Y=3080 $dt=1
M9 10 B 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3910 $Y=3080 $dt=1
M10 VDD 6 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4630 $Y=3080 $dt=1
M11 7 B VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5470 $Y=3080 $dt=1
.ends XNOR2X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OAI31XL                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OAI31XL A0 VDD VSS A1 A2 B0 Y
** N=10 EP=7 FDC=8
M0 8 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=760 $Y=1050 $dt=0
M1 VSS A1 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1600 $Y=1050 $dt=0
M2 8 A2 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2440 $Y=1050 $dt=0
M3 Y B0 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3280 $Y=1050 $dt=0
M4 9 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1360 $Y=3450 $dt=1
M5 10 A1 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1800 $Y=3450 $dt=1
M6 Y A2 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2440 $Y=3450 $dt=1
M7 VDD B0 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3280 $Y=3450 $dt=1
.ends OAI31XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AOI31XL                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AOI31XL A1 A0 VDD VSS A2 B0 Y
** N=10 EP=7 FDC=8
M0 8 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=880 $Y=1050 $dt=0
M1 9 A1 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1670 $Y=1050 $dt=0
M2 Y A2 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2350 $Y=1050 $dt=0
M3 VSS B0 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3190 $Y=1050 $dt=0
M4 10 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=830 $Y=2890 $dt=1
M5 VDD A1 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1670 $Y=2890 $dt=1
M6 10 A2 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2750 $Y=2890 $dt=1
M7 Y B0 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3590 $Y=2890 $dt=1
.ends AOI31XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AOI211XL                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AOI211XL A0 A1 VDD VSS Y B0 C0
** N=10 EP=7 FDC=8
M0 8 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1030 $dt=0
M1 Y A1 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1150 $Y=1030 $dt=0
M2 VSS B0 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1990 $Y=1030 $dt=0
M3 Y C0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2830 $Y=1030 $dt=0
M4 VDD A0 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=3380 $dt=1
M5 9 A1 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=3380 $dt=1
M6 10 B0 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2390 $Y=3380 $dt=1
M7 Y C0 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2830 $Y=3380 $dt=1
.ends AOI211XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AOI32XL                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AOI32XL A0 VDD VSS A1 A2 Y B1 B0
** N=12 EP=8 FDC=10
M0 9 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=880 $Y=830 $dt=0
M1 10 A1 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1520 $Y=830 $dt=0
M2 Y A2 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2240 $Y=830 $dt=0
M3 11 B1 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3470 $Y=830 $dt=0
M4 VSS B0 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3910 $Y=830 $dt=0
M5 12 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=830 $Y=2870 $dt=1
M6 VDD A1 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1670 $Y=2870 $dt=1
M7 12 A2 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2630 $Y=2870 $dt=1
M8 Y B1 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3470 $Y=2870 $dt=1
M9 12 B0 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4310 $Y=2870 $dt=1
.ends AOI32XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ACHCONX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ACHCONX2 A VDD VSS B CON CI
** N=13 EP=6 FDC=44
M0 10 A VSS VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=860 $Y=800 $dt=0
M1 VSS A 10 VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=1940 $Y=800 $dt=0
M2 11 10 VSS VSS nmos1v L=1e-07 W=2.6e-07 fw=2.6e-07 simw=2.6e-07 $X=3020 $Y=800 $dt=0
M3 VSS 10 11 VSS nmos1v L=1e-07 W=2.6e-07 fw=2.6e-07 simw=2.6e-07 $X=4100 $Y=800 $dt=0
M4 9 B VSS VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=5180 $Y=800 $dt=0
M5 VSS B 9 VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=6260 $Y=800 $dt=0
M6 8 9 10 VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=8120 $Y=800 $dt=0
M7 10 9 8 VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=9200 $Y=800 $dt=0
M8 7 B 10 VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=10280 $Y=800 $dt=0
M9 10 B 7 VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=11360 $Y=800 $dt=0
M10 7 9 11 VSS nmos1v L=1e-07 W=2.6e-07 fw=2.6e-07 simw=2.6e-07 $X=13220 $Y=840 $dt=0
M11 11 9 7 VSS nmos1v L=1e-07 W=2.6e-07 fw=2.6e-07 simw=2.6e-07 $X=14300 $Y=840 $dt=0
M12 8 B 11 VSS nmos1v L=1e-07 W=2.6e-07 fw=2.6e-07 simw=2.6e-07 $X=15860 $Y=840 $dt=0
M13 11 B 8 VSS nmos1v L=1e-07 W=2.6e-07 fw=2.6e-07 simw=2.6e-07 $X=16940 $Y=840 $dt=0
M14 12 B VSS VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=18800 $Y=800 $dt=0
M15 VSS B 12 VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=19880 $Y=800 $dt=0
M16 12 8 CON VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=21740 $Y=800 $dt=0
M17 CON 8 12 VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=22820 $Y=800 $dt=0
M18 13 7 CON VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=23900 $Y=800 $dt=0
M19 CON 7 13 VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=24980 $Y=800 $dt=0
M20 13 CI VSS VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=26840 $Y=800 $dt=0
M21 VSS CI 13 VSS nmos1v L=1e-07 W=3.25e-07 fw=3.25e-07 simw=3.25e-07 $X=27920 $Y=800 $dt=0
M22 10 A VDD VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=860 $Y=3130 $dt=1
M23 VDD A 10 VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=1940 $Y=3130 $dt=1
M24 11 10 VDD VDD pmos1v L=1e-07 W=4.3e-07 fw=4.3e-13 simw=4.3e-07 $X=3020 $Y=3560 $dt=1
M25 VDD 10 11 VDD pmos1v L=1e-07 W=4.3e-07 fw=4.3e-13 simw=4.3e-07 $X=4100 $Y=3560 $dt=1
M26 9 B VDD VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=5180 $Y=3130 $dt=1
M27 VDD B 9 VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=6260 $Y=3130 $dt=1
M28 8 B 10 VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=8120 $Y=3130 $dt=1
M29 10 B 8 VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=9200 $Y=3130 $dt=1
M30 7 9 10 VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=10280 $Y=3130 $dt=1
M31 10 9 7 VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=11360 $Y=3130 $dt=1
M32 7 B 11 VDD pmos1v L=1e-07 W=4.3e-07 fw=4.3e-13 simw=4.3e-07 $X=13220 $Y=3560 $dt=1
M33 11 B 7 VDD pmos1v L=1e-07 W=4.3e-07 fw=4.3e-13 simw=4.3e-07 $X=14300 $Y=3560 $dt=1
M34 8 9 11 VDD pmos1v L=1e-07 W=4.3e-07 fw=4.3e-13 simw=4.3e-07 $X=15860 $Y=3560 $dt=1
M35 11 9 8 VDD pmos1v L=1e-07 W=4.3e-07 fw=4.3e-13 simw=4.3e-07 $X=16940 $Y=3560 $dt=1
M36 12 B VDD VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=18800 $Y=3130 $dt=1
M37 VDD B 12 VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=19880 $Y=3130 $dt=1
M38 12 7 CON VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=21740 $Y=3130 $dt=1
M39 CON 7 12 VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=22820 $Y=3130 $dt=1
M40 13 8 CON VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=23900 $Y=3130 $dt=1
M41 CON 8 13 VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=24980 $Y=3130 $dt=1
M42 13 CI VDD VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=26840 $Y=3130 $dt=1
M43 VDD CI 13 VDD pmos1v L=1e-07 W=6.45e-07 fw=6.45e-13 simw=6.45e-07 $X=27920 $Y=3130 $dt=1
.ends ACHCONX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND4XL                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND4XL D VDD VSS C B A Y
** N=11 EP=7 FDC=10
M0 9 D 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1110 $Y=990 $dt=0
M1 10 C 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1550 $Y=990 $dt=0
M2 11 B 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2190 $Y=990 $dt=0
M3 VSS A 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2630 $Y=990 $dt=0
M4 Y 8 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3470 $Y=990 $dt=0
M5 8 D VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=3180 $dt=1
M6 VDD C 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=3180 $dt=1
M7 8 B VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2390 $Y=3180 $dt=1
M8 VDD A 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3230 $Y=3180 $dt=1
M9 Y 8 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4310 $Y=3180 $dt=1
.ends AND4XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR4XL                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR4XL D C VDD VSS B A Y
** N=11 EP=7 FDC=10
M0 8 D VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=720 $Y=1320 $dt=0
M1 VSS C 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1560 $Y=1320 $dt=0
M2 8 B VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2560 $Y=1320 $dt=0
M3 VSS A 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3400 $Y=1320 $dt=0
M4 Y 8 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4240 $Y=1320 $dt=0
M5 9 D 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=880 $Y=3440 $dt=1
M6 10 C 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1560 $Y=3440 $dt=1
M7 11 B 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2520 $Y=3440 $dt=1
M8 VDD A 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2960 $Y=3440 $dt=1
M9 Y 8 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3800 $Y=3440 $dt=1
.ends OR4XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO22X1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO22X1 A0 VDD VSS A1 B1 B0 Y
** N=11 EP=7 FDC=10
M0 9 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1310 $Y=1180 $dt=0
M1 8 A1 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1750 $Y=1180 $dt=0
M2 10 B1 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2590 $Y=1180 $dt=0
M3 VSS B0 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3390 $Y=1180 $dt=0
M4 Y 8 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=4350 $Y=800 $dt=0
M5 VDD A0 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=2880 $dt=1
M6 11 A1 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1750 $Y=2880 $dt=1
M7 8 B1 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2590 $Y=2880 $dt=1
M8 11 B0 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3430 $Y=2880 $dt=1
M9 Y 8 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=4890 $Y=3120 $dt=1
.ends AO22X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND4X1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND4X1 D C VDD VSS B A Y
** N=11 EP=7 FDC=10
M0 9 D 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=880 $Y=1220 $dt=0
M1 10 C 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1520 $Y=1220 $dt=0
M2 11 B 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2630 $Y=1220 $dt=0
M3 VSS A 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3070 $Y=1220 $dt=0
M4 Y 8 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=4030 $Y=840 $dt=0
M5 8 D VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=3000 $dt=1
M6 VDD C 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=3000 $dt=1
M7 8 B VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2630 $Y=3000 $dt=1
M8 VDD A 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3470 $Y=3000 $dt=1
M9 Y 8 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=4310 $Y=2680 $dt=1
.ends AND4X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR4X1                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR4X1 D C VDD VSS B A Y
** N=11 EP=7 FDC=10
M0 8 D VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1320 $dt=0
M1 VSS C 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1550 $Y=1320 $dt=0
M2 8 B VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2510 $Y=1320 $dt=0
M3 VSS A 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3350 $Y=1320 $dt=0
M4 Y 8 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=4310 $Y=940 $dt=0
M5 9 D 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1390 $Y=3160 $dt=1
M6 10 C 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1830 $Y=3160 $dt=1
M7 11 B 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2510 $Y=3160 $dt=1
M8 VDD A 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3350 $Y=3160 $dt=1
M9 Y 8 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=4310 $Y=3120 $dt=1
.ends OR4X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OAI222XL                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OAI222XL A0 A1 VDD VSS B0 B1 C0 Y C1
** N=14 EP=9 FDC=12
M0 10 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=610 $Y=1320 $dt=0
M1 VSS A1 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1450 $Y=1320 $dt=0
M2 10 B1 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2950 $Y=1200 $dt=0
M3 11 B0 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3790 $Y=1200 $dt=0
M4 Y C0 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4630 $Y=1200 $dt=0
M5 11 C1 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5470 $Y=1200 $dt=0
M6 12 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1010 $Y=3700 $dt=1
M7 Y A1 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1450 $Y=3700 $dt=1
M8 13 B1 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2950 $Y=3700 $dt=1
M9 VDD B0 13 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3790 $Y=3700 $dt=1
M10 14 C0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4630 $Y=3700 $dt=1
M11 Y C1 14 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5070 $Y=3700 $dt=1
.ends OAI222XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OA22X1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OA22X1 A0 A1 VDD VSS B1 B0 Y
** N=11 EP=7 FDC=10
M0 VSS A0 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1360 $dt=0
M1 9 A1 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1710 $Y=1360 $dt=0
M2 8 B1 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2550 $Y=1360 $dt=0
M3 9 B0 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3390 $Y=1360 $dt=0
M4 Y 8 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=4890 $Y=800 $dt=0
M5 10 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=880 $Y=3240 $dt=1
M6 8 A1 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1710 $Y=3240 $dt=1
M7 11 B1 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2550 $Y=3240 $dt=1
M8 VDD B0 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3190 $Y=3240 $dt=1
M9 Y 8 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=4150 $Y=3120 $dt=1
.ends OA22X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2BX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2BX1 Y B VDD VSS AN
** N=7 EP=5 FDC=6
M0 7 B Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1120 $Y=800 $dt=0
M1 VSS 6 7 VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1560 $Y=800 $dt=0
M2 6 AN VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2520 $Y=1180 $dt=0
M3 Y B VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=840 $Y=3120 $dt=1
M4 VDD 6 Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1680 $Y=3120 $dt=1
M5 6 AN VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2520 $Y=3240 $dt=1
.ends NAND2BX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MX2X1                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MX2X1 S0 A VDD VSS B Y
** N=12 EP=6 FDC=12
M0 VSS S0 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=800 $dt=0
M1 9 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1550 $Y=800 $dt=0
M2 7 8 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1990 $Y=800 $dt=0
M3 10 S0 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2830 $Y=800 $dt=0
M4 VSS B 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3270 $Y=800 $dt=0
M5 Y 7 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=4110 $Y=800 $dt=0
M6 VDD S0 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=3600 $dt=1
M7 11 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=3600 $dt=1
M8 7 S0 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1990 $Y=3600 $dt=1
M9 12 8 7 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2830 $Y=3600 $dt=1
M10 VDD B 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3270 $Y=3600 $dt=1
M11 Y 7 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=4230 $Y=3120 $dt=1
.ends MX2X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AOI2BB1X1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AOI2BB1X1 Y VDD VSS B0 A0N A1N
** N=9 EP=6 FDC=8
M0 Y 7 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=920 $Y=880 $dt=0
M1 VSS B0 Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1760 $Y=880 $dt=0
M2 7 A0N VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2600 $Y=1240 $dt=0
M3 VSS A1N 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3440 $Y=1240 $dt=0
M4 8 7 Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1200 $Y=3120 $dt=1
M5 VDD B0 8 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1640 $Y=3120 $dt=1
M6 9 A0N VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2600 $Y=3120 $dt=1
M7 7 A1N 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3040 $Y=3120 $dt=1
.ends AOI2BB1X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OAI2BB1X1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OAI2BB1X1 Y VDD VSS B0 A0N A1N
** N=9 EP=6 FDC=8
M0 8 7 Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=950 $Y=820 $dt=0
M1 VSS B0 8 VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1550 $Y=820 $dt=0
M2 9 A0N VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2510 $Y=1200 $dt=0
M3 7 A1N 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2980 $Y=1200 $dt=0
M4 Y 7 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=3080 $dt=1
M5 VDD B0 Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1550 $Y=3080 $dt=1
M6 7 A0N VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2390 $Y=3180 $dt=1
M7 VDD A1N 7 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3230 $Y=3180 $dt=1
.ends OAI2BB1X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NOR2XL                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NOR2XL A B Y VDD VSS
** N=6 EP=5 FDC=4
M0 Y A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=590 $Y=1330 $dt=0
M1 VSS B Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1430 $Y=1330 $dt=0
M2 6 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=750 $Y=3170 $dt=1
M3 Y B 6 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1190 $Y=3170 $dt=1
.ends NOR2XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INVXL                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INVXL A Y VDD VSS
** N=4 EP=4 FDC=2
M0 Y A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1360 $dt=0
M1 Y A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=2910 $dt=1
.ends INVXL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NOR4BBX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NOR4BBX1 BN VDD VSS D Y C AN
** N=12 EP=7 FDC=12
M0 9 BN VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=650 $Y=1360 $dt=0
M1 Y D VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=2110 $Y=800 $dt=0
M2 VSS C Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=2950 $Y=800 $dt=0
M3 Y 9 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=3790 $Y=800 $dt=0
M4 VSS 8 Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=4630 $Y=800 $dt=0
M5 8 AN VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5470 $Y=1180 $dt=0
M6 9 BN VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=720 $Y=2680 $dt=1
M7 10 D Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=2340 $Y=3120 $dt=1
M8 11 C 10 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=2950 $Y=3120 $dt=1
M9 12 9 11 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=3420 $Y=3120 $dt=1
M10 VDD 8 12 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=3860 $Y=3120 $dt=1
M11 8 AN VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5300 $Y=3120 $dt=1
.ends NOR4BBX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND2X1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND2X1 B VDD VSS A Y
** N=7 EP=5 FDC=6
M0 7 B 6 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=830 $Y=1220 $dt=0
M1 VSS A 7 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1270 $Y=1220 $dt=0
M2 Y 6 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=2230 $Y=840 $dt=0
M3 6 B VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=3250 $dt=1
M4 VDD A 6 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=3250 $dt=1
M5 Y 6 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=2390 $Y=2680 $dt=1
.ends AND2X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__P1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__P1 1 2 3 4 12 13 14 15 16 17
+ 18 19 20 21 22 23 24 25 26 27
+ 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47
+ 48 49 50 51 52 53 55 56 57 58
+ 59 60 61 62 63 64 65 66 67 68
+ 69 70 71 72 73 74 75 76 77 78
+ 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 96 97 98 99
+ 100 101 102 103 104 106 107 108 109 110
+ 111 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 127 128 129 130 131 132
+ 134 135 136 137 138 140 141 142 143 144
+ 145 146 148 149 150 151 152 153 154 155
+ 156 158 159 160 161 162 163 164 165 167
+ 168 169 170 172 173 174 176 177 178 179
+ 180 181 183 184 185 186 187 188 189 190
+ 191 192 193 194 196 197 198 199
** N=1663 EP=178 FDC=21518
X0 207 13 12 2 CLKBUFX2 $T=34800 157180 1 0 $X=34200 $Y=151360
X1 208 13 12 19 CLKBUFX2 $T=35380 52780 1 0 $X=34780 $Y=46960
X2 209 13 12 4 CLKBUFX2 $T=35960 63220 1 0 $X=35360 $Y=57400
X3 210 13 12 16 CLKBUFX2 $T=35960 84100 0 0 $X=35360 $Y=83740
X4 211 13 12 3 CLKBUFX2 $T=36540 146740 1 0 $X=35940 $Y=140920
X5 212 13 12 18 CLKBUFX2 $T=37120 115420 1 0 $X=36520 $Y=109600
X6 213 13 12 1 CLKBUFX2 $T=37120 136300 1 0 $X=36520 $Y=130480
X7 214 13 12 15 CLKBUFX2 $T=37700 115420 0 0 $X=37100 $Y=115060
X8 215 13 12 21 CLKBUFX2 $T=38280 21460 1 0 $X=37680 $Y=15640
X9 216 13 12 20 CLKBUFX2 $T=38860 31900 0 0 $X=38260 $Y=31540
X10 217 13 12 14 CLKBUFX2 $T=39440 73660 0 0 $X=38840 $Y=73300
X11 218 13 12 17 CLKBUFX2 $T=40600 136300 1 0 $X=40000 $Y=130480
X12 219 13 12 27 CLKBUFX2 $T=48720 21460 1 0 $X=48120 $Y=15640
X13 220 13 12 25 CLKBUFX2 $T=55100 31900 1 0 $X=54500 $Y=26080
X14 221 13 12 51 CLKBUFX2 $T=110780 21460 0 0 $X=110180 $Y=21100
X15 222 13 12 75 CLKBUFX2 $T=176320 31900 1 0 $X=175720 $Y=26080
X16 70 13 12 24 CLKINVX2 $T=164720 115420 1 0 $X=164120 $Y=109600
X17 70 13 12 118 CLKINVX2 $T=370620 63220 1 180 $X=367120 $Y=62860
X18 199 13 12 141 CLKINVX2 $T=546360 21460 0 180 $X=542860 $Y=15640
X19 223 224 13 12 CLKINVX1 $T=49300 115420 0 0 $X=48700 $Y=115060
X20 225 226 13 12 CLKINVX1 $T=58000 146740 1 0 $X=57400 $Y=140920
X21 227 228 13 12 CLKINVX1 $T=58580 115420 1 0 $X=57980 $Y=109600
X22 229 230 13 12 CLKINVX1 $T=59740 52780 1 0 $X=59140 $Y=46960
X23 32 231 13 12 CLKINVX1 $T=64380 167620 1 180 $X=62040 $Y=167260
X24 232 233 13 12 CLKINVX1 $T=68440 136300 1 180 $X=66100 $Y=135940
X25 234 235 13 12 CLKINVX1 $T=67860 125860 1 0 $X=67260 $Y=120040
X26 236 237 13 12 CLKINVX1 $T=68440 42340 0 0 $X=67840 $Y=41980
X27 238 239 13 12 CLKINVX1 $T=71920 63220 1 0 $X=71320 $Y=57400
X28 240 241 13 12 CLKINVX1 $T=73660 73660 0 0 $X=73060 $Y=73300
X29 242 243 13 12 CLKINVX1 $T=74240 167620 0 0 $X=73640 $Y=167260
X30 244 245 13 12 CLKINVX1 $T=81780 73660 0 180 $X=79440 $Y=67840
X31 246 247 13 12 CLKINVX1 $T=85840 104980 0 180 $X=83500 $Y=99160
X32 248 37 13 12 CLKINVX1 $T=85840 178060 1 180 $X=83500 $Y=177700
X33 249 250 13 12 CLKINVX1 $T=86420 125860 0 180 $X=84080 $Y=120040
X34 251 252 13 12 CLKINVX1 $T=91640 63220 0 180 $X=89300 $Y=57400
X35 253 254 13 12 CLKINVX1 $T=91060 94540 1 0 $X=90460 $Y=88720
X36 255 256 13 12 CLKINVX1 $T=100920 73660 0 0 $X=100320 $Y=73300
X37 46 257 13 12 CLKINVX1 $T=105560 178060 0 180 $X=103220 $Y=172240
X38 258 259 13 12 CLKINVX1 $T=111360 73660 1 0 $X=110760 $Y=67840
X39 260 261 13 12 CLKINVX1 $T=113100 104980 0 180 $X=110760 $Y=99160
X40 262 263 13 12 CLKINVX1 $T=116580 73660 0 180 $X=114240 $Y=67840
X41 264 265 13 12 CLKINVX1 $T=118320 115420 0 180 $X=115980 $Y=109600
X42 55 266 13 12 CLKINVX1 $T=125860 157180 0 0 $X=125260 $Y=156820
X43 267 268 13 12 CLKINVX1 $T=128180 42340 0 180 $X=125840 $Y=36520
X44 269 270 13 12 CLKINVX1 $T=126440 178060 0 0 $X=125840 $Y=177700
X45 271 272 13 12 CLKINVX1 $T=127600 52780 0 0 $X=127000 $Y=52420
X46 273 274 13 12 CLKINVX1 $T=128760 125860 1 0 $X=128160 $Y=120040
X47 57 275 13 12 CLKINVX1 $T=134560 188500 0 180 $X=132220 $Y=182680
X48 276 277 13 12 CLKINVX1 $T=133400 31900 1 0 $X=132800 $Y=26080
X49 278 279 13 12 CLKINVX1 $T=133400 157180 0 0 $X=132800 $Y=156820
X50 280 281 13 12 CLKINVX1 $T=133400 178060 0 0 $X=132800 $Y=177700
X51 282 283 13 12 CLKINVX1 $T=138040 178060 1 0 $X=137440 $Y=172240
X52 284 61 13 12 CLKINVX1 $T=142680 188500 1 0 $X=142080 $Y=182680
X53 285 286 13 12 CLKINVX1 $T=145000 104980 1 180 $X=142660 $Y=104620
X54 287 288 13 12 CLKINVX1 $T=145580 73660 1 0 $X=144980 $Y=67840
X55 289 290 13 12 CLKINVX1 $T=145580 178060 0 0 $X=144980 $Y=177700
X56 291 292 13 12 CLKINVX1 $T=146740 157180 1 0 $X=146140 $Y=151360
X57 293 294 13 12 CLKINVX1 $T=147900 63220 1 0 $X=147300 $Y=57400
X58 295 296 13 12 CLKINVX1 $T=149640 178060 1 180 $X=147300 $Y=177700
X59 297 298 13 12 CLKINVX1 $T=149640 136300 1 0 $X=149040 $Y=130480
X60 299 300 13 12 CLKINVX1 $T=150800 52780 0 0 $X=150200 $Y=52420
X61 301 302 13 12 CLKINVX1 $T=158340 94540 1 180 $X=156000 $Y=94180
X62 303 304 13 12 CLKINVX1 $T=156600 167620 1 0 $X=156000 $Y=161800
X63 305 306 13 12 CLKINVX1 $T=157760 167620 0 0 $X=157160 $Y=167260
X64 307 308 13 12 CLKINVX1 $T=158340 104980 1 0 $X=157740 $Y=99160
X65 309 310 13 12 CLKINVX1 $T=158340 167620 1 0 $X=157740 $Y=161800
X66 311 312 13 12 CLKINVX1 $T=158920 146740 0 0 $X=158320 $Y=146380
X67 313 314 13 12 CLKINVX1 $T=161240 157180 0 0 $X=160640 $Y=156820
X68 70 315 13 12 CLKINVX1 $T=162980 115420 1 0 $X=162380 $Y=109600
X69 316 317 13 12 CLKINVX1 $T=166460 52780 1 180 $X=164120 $Y=52420
X70 318 319 13 12 CLKINVX1 $T=173420 104980 0 0 $X=172820 $Y=104620
X71 70 320 13 12 CLKINVX1 $T=174000 115420 1 0 $X=173400 $Y=109600
X72 76 321 13 12 CLKINVX1 $T=177480 167620 1 0 $X=176880 $Y=161800
X73 322 323 13 12 CLKINVX1 $T=179800 136300 1 0 $X=179200 $Y=130480
X74 324 325 13 12 CLKINVX1 $T=186180 84100 0 0 $X=185580 $Y=83740
X75 326 327 13 12 CLKINVX1 $T=188500 84100 0 180 $X=186160 $Y=78280
X76 328 329 13 12 CLKINVX1 $T=191400 63220 0 180 $X=189060 $Y=57400
X77 81 330 13 12 CLKINVX1 $T=194300 178060 0 180 $X=191960 $Y=172240
X78 331 332 13 12 CLKINVX1 $T=194880 73660 1 180 $X=192540 $Y=73300
X79 333 334 13 12 CLKINVX1 $T=193140 146740 0 0 $X=192540 $Y=146380
X80 335 336 13 12 CLKINVX1 $T=200100 63220 0 180 $X=197760 $Y=57400
X81 337 338 13 12 CLKINVX1 $T=198360 94540 0 0 $X=197760 $Y=94180
X82 339 340 13 12 CLKINVX1 $T=201260 42340 1 180 $X=198920 $Y=41980
X83 341 342 13 12 CLKINVX1 $T=201260 157180 0 180 $X=198920 $Y=151360
X84 84 343 13 12 CLKINVX1 $T=200680 167620 1 0 $X=200080 $Y=161800
X85 344 345 13 12 CLKINVX1 $T=206480 73660 0 0 $X=205880 $Y=73300
X86 346 347 13 12 CLKINVX1 $T=207640 52780 1 0 $X=207040 $Y=46960
X87 70 85 13 12 CLKINVX1 $T=210540 115420 1 0 $X=209940 $Y=109600
X88 348 349 13 12 CLKINVX1 $T=215180 31900 1 180 $X=212840 $Y=31540
X89 86 350 13 12 CLKINVX1 $T=216920 178060 1 180 $X=214580 $Y=177700
X90 351 352 13 12 CLKINVX1 $T=223880 115420 0 180 $X=221540 $Y=109600
X91 353 354 13 12 CLKINVX1 $T=222720 136300 1 0 $X=222120 $Y=130480
X92 355 356 13 12 CLKINVX1 $T=225040 167620 1 0 $X=224440 $Y=161800
X93 357 358 13 12 CLKINVX1 $T=229100 104980 1 180 $X=226760 $Y=104620
X94 359 360 13 12 CLKINVX1 $T=229100 115420 0 180 $X=226760 $Y=109600
X95 361 362 13 12 CLKINVX1 $T=227360 136300 0 0 $X=226760 $Y=135940
X96 363 364 13 12 CLKINVX1 $T=227940 167620 1 0 $X=227340 $Y=161800
X97 365 366 13 12 CLKINVX1 $T=230840 125860 1 0 $X=230240 $Y=120040
X98 367 368 13 12 CLKINVX1 $T=230840 167620 1 0 $X=230240 $Y=161800
X99 369 370 13 12 CLKINVX1 $T=232580 73660 1 0 $X=231980 $Y=67840
X100 371 372 13 12 CLKINVX1 $T=234320 125860 0 0 $X=233720 $Y=125500
X101 373 374 13 12 CLKINVX1 $T=236060 136300 1 180 $X=233720 $Y=135940
X102 375 376 13 12 CLKINVX1 $T=234900 21460 0 0 $X=234300 $Y=21100
X103 377 378 13 12 CLKINVX1 $T=240120 115420 1 0 $X=239520 $Y=109600
X104 379 380 13 12 CLKINVX1 $T=243020 115420 1 180 $X=240680 $Y=115060
X105 381 382 13 12 CLKINVX1 $T=243020 104980 1 0 $X=242420 $Y=99160
X106 383 384 13 12 CLKINVX1 $T=245340 125860 0 0 $X=244740 $Y=125500
X107 385 386 13 12 CLKINVX1 $T=246500 52780 1 0 $X=245900 $Y=46960
X108 387 388 13 12 CLKINVX1 $T=248820 42340 0 180 $X=246480 $Y=36520
X109 389 390 13 12 CLKINVX1 $T=254040 125860 1 0 $X=253440 $Y=120040
X110 391 392 13 12 CLKINVX1 $T=256940 52780 1 0 $X=256340 $Y=46960
X111 393 394 13 12 CLKINVX1 $T=258100 21460 1 0 $X=257500 $Y=15640
X112 395 396 13 12 CLKINVX1 $T=258100 31900 0 0 $X=257500 $Y=31540
X113 397 398 13 12 CLKINVX1 $T=260420 52780 1 0 $X=259820 $Y=46960
X114 399 400 13 12 CLKINVX1 $T=262160 125860 0 180 $X=259820 $Y=120040
X115 401 402 13 12 CLKINVX1 $T=261580 73660 1 0 $X=260980 $Y=67840
X116 403 404 13 12 CLKINVX1 $T=263320 94540 1 180 $X=260980 $Y=94180
X117 405 406 13 12 CLKINVX1 $T=265640 31900 1 0 $X=265040 $Y=26080
X118 407 408 13 12 CLKINVX1 $T=271440 42340 0 0 $X=270840 $Y=41980
X119 110 409 13 12 CLKINVX1 $T=277240 178060 1 180 $X=274900 $Y=177700
X120 410 411 13 12 CLKINVX1 $T=278400 157180 0 180 $X=276060 $Y=151360
X121 412 413 13 12 CLKINVX1 $T=280720 167620 0 0 $X=280120 $Y=167260
X122 414 415 13 12 CLKINVX1 $T=283040 104980 0 180 $X=280700 $Y=99160
X123 416 417 13 12 CLKINVX1 $T=288260 84100 1 0 $X=287660 $Y=78280
X124 418 419 13 12 CLKINVX1 $T=290000 73660 1 0 $X=289400 $Y=67840
X125 420 421 13 12 CLKINVX1 $T=294060 136300 1 180 $X=291720 $Y=135940
X126 422 423 13 12 CLKINVX1 $T=296960 115420 0 180 $X=294620 $Y=109600
X127 424 425 13 12 CLKINVX1 $T=295800 104980 1 0 $X=295200 $Y=99160
X128 426 427 13 12 CLKINVX1 $T=302760 188500 1 0 $X=302160 $Y=182680
X129 428 429 13 12 CLKINVX1 $T=305080 42340 1 0 $X=304480 $Y=36520
X130 430 431 13 12 CLKINVX1 $T=305080 115420 0 0 $X=304480 $Y=115060
X131 432 433 13 12 CLKINVX1 $T=309720 73660 0 180 $X=307380 $Y=67840
X132 434 435 13 12 CLKINVX1 $T=310880 52780 1 0 $X=310280 $Y=46960
X133 436 437 13 12 CLKINVX1 $T=313200 42340 0 180 $X=310860 $Y=36520
X134 438 439 13 12 CLKINVX1 $T=316100 73660 1 0 $X=315500 $Y=67840
X135 440 441 13 12 CLKINVX1 $T=318420 146740 0 0 $X=317820 $Y=146380
X136 442 443 13 12 CLKINVX1 $T=319000 31900 1 0 $X=318400 $Y=26080
X137 444 445 13 12 CLKINVX1 $T=320160 42340 0 0 $X=319560 $Y=41980
X138 446 447 13 12 CLKINVX1 $T=321320 73660 1 0 $X=320720 $Y=67840
X139 448 449 13 12 CLKINVX1 $T=329440 104980 0 180 $X=327100 $Y=99160
X140 450 451 13 12 CLKINVX1 $T=340460 104980 0 180 $X=338120 $Y=99160
X141 452 453 13 12 CLKINVX1 $T=345680 178060 1 180 $X=343340 $Y=177700
X142 454 455 13 12 CLKINVX1 $T=346840 84100 0 0 $X=346240 $Y=83740
X143 456 457 13 12 CLKINVX1 $T=346840 178060 0 0 $X=346240 $Y=177700
X144 458 459 13 12 CLKINVX1 $T=357280 73660 0 0 $X=356680 $Y=73300
X145 460 461 13 12 CLKINVX1 $T=360760 63220 0 180 $X=358420 $Y=57400
X146 462 463 13 12 CLKINVX1 $T=361920 42340 1 0 $X=361320 $Y=36520
X147 464 465 13 12 CLKINVX1 $T=363660 42340 1 0 $X=363060 $Y=36520
X148 466 467 13 12 CLKINVX1 $T=364820 21460 0 0 $X=364220 $Y=21100
X149 468 469 13 12 CLKINVX1 $T=370040 42340 0 0 $X=369440 $Y=41980
X150 470 471 13 12 CLKINVX1 $T=372940 94540 1 180 $X=370600 $Y=94180
X151 472 473 13 12 CLKINVX1 $T=378740 178060 0 0 $X=378140 $Y=177700
X152 70 474 13 12 CLKINVX1 $T=379320 73660 1 0 $X=378720 $Y=67840
X153 475 476 13 12 CLKINVX1 $T=379320 73660 0 0 $X=378720 $Y=73300
X154 477 478 13 12 CLKINVX1 $T=379320 94540 0 0 $X=378720 $Y=94180
X155 479 480 13 12 CLKINVX1 $T=379900 125860 0 0 $X=379300 $Y=125500
X156 141 70 13 12 CLKINVX1 $T=381060 63220 0 0 $X=380460 $Y=62860
X157 481 482 13 12 CLKINVX1 $T=381640 136300 0 0 $X=381040 $Y=135940
X158 483 484 13 12 CLKINVX1 $T=381640 157180 1 0 $X=381040 $Y=151360
X159 485 486 13 12 CLKINVX1 $T=385700 104980 1 180 $X=383360 $Y=104620
X160 487 488 13 12 CLKINVX1 $T=388600 136300 0 180 $X=386260 $Y=130480
X161 489 490 13 12 CLKINVX1 $T=387440 125860 1 0 $X=386840 $Y=120040
X162 491 492 13 12 CLKINVX1 $T=388020 115420 1 0 $X=387420 $Y=109600
X163 493 494 13 12 CLKINVX1 $T=391500 42340 1 180 $X=389160 $Y=41980
X164 495 496 13 12 CLKINVX1 $T=393820 125860 0 0 $X=393220 $Y=125500
X165 497 498 13 12 CLKINVX1 $T=395560 188500 1 0 $X=394960 $Y=182680
X166 499 500 13 12 CLKINVX1 $T=397880 125860 1 180 $X=395540 $Y=125500
X167 501 502 13 12 CLKINVX1 $T=399040 115420 1 0 $X=398440 $Y=109600
X168 503 504 13 12 CLKINVX1 $T=399040 125860 0 0 $X=398440 $Y=125500
X169 505 506 13 12 CLKINVX1 $T=400780 115420 1 0 $X=400180 $Y=109600
X170 507 508 13 12 CLKINVX1 $T=403680 84100 1 180 $X=401340 $Y=83740
X171 509 510 13 12 CLKINVX1 $T=405420 52780 1 0 $X=404820 $Y=46960
X172 511 512 13 12 CLKINVX1 $T=407160 136300 1 0 $X=406560 $Y=130480
X173 513 514 13 12 CLKINVX1 $T=408320 63220 1 0 $X=407720 $Y=57400
X174 515 516 13 12 CLKINVX1 $T=408900 125860 0 0 $X=408300 $Y=125500
X175 517 518 13 12 CLKINVX1 $T=411800 84100 0 180 $X=409460 $Y=78280
X176 519 520 13 12 CLKINVX1 $T=416440 104980 0 0 $X=415840 $Y=104620
X177 521 522 13 12 CLKINVX1 $T=417600 115420 1 0 $X=417000 $Y=109600
X178 523 524 13 12 CLKINVX1 $T=420500 157180 1 180 $X=418160 $Y=156820
X179 525 526 13 12 CLKINVX1 $T=419340 94540 0 0 $X=418740 $Y=94180
X180 527 528 13 12 CLKINVX1 $T=430360 157180 1 180 $X=428020 $Y=156820
X181 529 530 13 12 CLKINVX1 $T=440800 52780 0 0 $X=440200 $Y=52420
X182 531 532 13 12 CLKINVX1 $T=441960 73660 1 0 $X=441360 $Y=67840
X183 533 534 13 12 CLKINVX1 $T=443700 84100 0 0 $X=443100 $Y=83740
X184 535 536 13 12 CLKINVX1 $T=444280 104980 1 0 $X=443680 $Y=99160
X185 537 538 13 12 CLKINVX1 $T=446020 136300 1 180 $X=443680 $Y=135940
X186 539 540 13 12 CLKINVX1 $T=446600 178060 0 180 $X=444260 $Y=172240
X187 541 160 13 12 CLKINVX1 $T=446600 188500 0 180 $X=444260 $Y=182680
X188 542 543 13 12 CLKINVX1 $T=447180 178060 1 0 $X=446580 $Y=172240
X189 544 545 13 12 CLKINVX1 $T=448920 94540 1 0 $X=448320 $Y=88720
X190 546 547 13 12 CLKINVX1 $T=449500 104980 1 0 $X=448900 $Y=99160
X191 548 549 13 12 CLKINVX1 $T=450080 31900 0 0 $X=449480 $Y=31540
X192 166 550 13 12 CLKINVX1 $T=453560 188500 0 180 $X=451220 $Y=182680
X193 551 552 13 12 CLKINVX1 $T=459940 178060 1 180 $X=457600 $Y=177700
X194 553 554 13 12 CLKINVX1 $T=459940 84100 0 0 $X=459340 $Y=83740
X195 555 556 13 12 CLKINVX1 $T=461680 104980 1 0 $X=461080 $Y=99160
X196 557 558 13 12 CLKINVX1 $T=469800 104980 1 180 $X=467460 $Y=104620
X197 559 560 13 12 CLKINVX1 $T=469220 178060 1 0 $X=468620 $Y=172240
X198 561 562 13 12 CLKINVX1 $T=472700 167620 0 0 $X=472100 $Y=167260
X199 563 564 13 12 CLKINVX1 $T=501120 42340 1 180 $X=498780 $Y=41980
X200 565 566 13 12 CLKINVX1 $T=501120 94540 1 0 $X=500520 $Y=88720
X201 567 568 13 12 CLKINVX1 $T=501700 31900 1 0 $X=501100 $Y=26080
X202 569 570 13 12 CLKINVX1 $T=504020 73660 0 180 $X=501680 $Y=67840
X203 571 572 13 12 CLKINVX1 $T=504020 21460 1 0 $X=503420 $Y=15640
X204 573 574 13 12 CLKINVX1 $T=504020 136300 1 0 $X=503420 $Y=130480
X205 575 576 13 12 CLKINVX1 $T=506920 115420 0 0 $X=506320 $Y=115060
X206 577 578 13 12 CLKINVX1 $T=507500 125860 0 0 $X=506900 $Y=125500
X207 579 580 13 12 CLKINVX1 $T=513300 136300 1 0 $X=512700 $Y=130480
X208 581 582 13 12 CLKINVX1 $T=515040 188500 1 0 $X=514440 $Y=182680
X209 583 584 13 12 CLKINVX1 $T=515620 125860 0 0 $X=515020 $Y=125500
X210 585 586 13 12 CLKINVX1 $T=517940 136300 0 180 $X=515600 $Y=130480
X211 587 588 13 12 CLKINVX1 $T=523160 178060 0 180 $X=520820 $Y=172240
X212 589 22 13 12 315 215 DFFRHQX1 $T=52200 21460 1 180 $X=35940 $Y=21100
X213 590 22 13 12 315 216 DFFRHQX1 $T=52780 31900 0 180 $X=36520 $Y=26080
X214 591 22 13 12 315 208 DFFRHQX1 $T=53360 42340 1 180 $X=37100 $Y=41980
X215 592 22 13 12 315 209 DFFRHQX1 $T=55100 63220 0 180 $X=38840 $Y=57400
X216 593 22 13 12 315 219 DFFRHQX1 $T=67860 21460 0 180 $X=51600 $Y=15640
X217 594 22 13 12 315 220 DFFRHQX1 $T=69020 21460 1 180 $X=52760 $Y=21100
X218 595 22 13 12 315 596 DFFRHQX1 $T=85840 31900 0 180 $X=69580 $Y=26080
X219 597 22 13 12 315 593 DFFRHQX1 $T=86420 21460 0 180 $X=70160 $Y=15640
X220 598 22 13 12 315 594 DFFRHQX1 $T=86420 21460 1 180 $X=70160 $Y=21100
X221 599 22 13 12 315 600 DFFRHQX1 $T=86420 42340 0 180 $X=70160 $Y=36520
X222 601 22 13 12 315 597 DFFRHQX1 $T=104980 21460 0 180 $X=88720 $Y=15640
X223 602 22 13 12 315 598 DFFRHQX1 $T=89900 21460 0 0 $X=89300 $Y=21100
X224 603 22 13 12 315 221 DFFRHQX1 $T=124700 21460 0 180 $X=108440 $Y=15640
X225 604 22 13 12 320 603 DFFRHQX1 $T=129920 21460 1 180 $X=113660 $Y=21100
X226 605 22 13 12 320 604 DFFRHQX1 $T=142100 21460 0 180 $X=125840 $Y=15640
X227 606 22 13 12 320 605 DFFRHQX1 $T=147900 21460 1 180 $X=131640 $Y=21100
X228 607 22 13 12 24 73 DFFRHQX1 $T=161820 136300 1 0 $X=161220 $Y=130480
X229 608 22 13 12 320 222 DFFRHQX1 $T=164140 21460 1 0 $X=163540 $Y=15640
X230 609 22 13 12 320 608 DFFRHQX1 $T=180380 21460 1 180 $X=164120 $Y=21100
X231 610 22 13 12 320 609 DFFRHQX1 $T=195460 31900 0 180 $X=179200 $Y=26080
X232 611 22 13 12 320 612 DFFRHQX1 $T=196040 21460 0 180 $X=179780 $Y=15640
X233 612 22 13 12 320 610 DFFRHQX1 $T=180380 21460 0 0 $X=179780 $Y=21100
X234 613 22 13 12 85 99 DFFRHQX1 $T=256940 178060 0 180 $X=240680 $Y=172240
X235 614 22 13 12 118 615 DFFRHQX1 $T=303920 31900 0 180 $X=287660 $Y=26080
X236 616 22 13 12 118 617 DFFRHQX1 $T=340460 73660 0 180 $X=324200 $Y=67840
X237 618 22 13 12 474 619 DFFRHQX1 $T=417600 21460 0 180 $X=401340 $Y=15640
X238 620 22 13 12 474 621 DFFRHQX1 $T=418180 21460 1 180 $X=401920 $Y=21100
X239 622 22 13 12 141 623 DFFRHQX1 $T=429780 157180 0 180 $X=413520 $Y=151360
X240 624 22 13 12 474 620 DFFRHQX1 $T=436740 21460 1 180 $X=420480 $Y=21100
X241 625 22 13 12 141 626 DFFRHQX1 $T=527220 21460 0 180 $X=510960 $Y=15640
X242 627 22 13 12 24 628 629 630 SDFFRHQX1 $T=105560 125860 1 180 $X=85820 $Y=125500
X243 631 22 13 12 85 345 344 632 SDFFRHQX1 $T=223880 84100 0 180 $X=204140 $Y=78280
X244 633 22 13 12 85 634 635 636 SDFFRHQX1 $T=279560 84100 1 180 $X=259820 $Y=83740
X245 637 13 12 638 22 315 210 DFFRX1 $T=51620 94540 0 180 $X=34200 $Y=88720
X246 639 13 12 640 22 24 218 DFFRX1 $T=51620 125860 1 180 $X=34200 $Y=125500
X247 641 13 12 642 22 315 212 DFFRX1 $T=52200 104980 0 180 $X=34780 $Y=99160
X248 643 13 12 644 22 24 213 DFFRX1 $T=52200 136300 1 180 $X=34780 $Y=135940
X249 645 13 12 646 22 24 214 DFFRX1 $T=52780 125860 0 180 $X=35360 $Y=120040
X250 647 13 12 648 22 315 589 DFFRX1 $T=54520 42340 0 180 $X=37100 $Y=36520
X251 649 13 12 650 22 315 217 DFFRX1 $T=54520 84100 0 180 $X=37100 $Y=78280
X252 651 13 12 652 22 24 211 DFFRX1 $T=54520 146740 1 180 $X=37100 $Y=146380
X253 653 13 12 23 22 24 207 DFFRX1 $T=55100 157180 0 180 $X=37680 $Y=151360
X254 654 13 12 655 22 315 591 DFFRX1 $T=55680 52780 0 180 $X=38260 $Y=46960
X255 656 13 12 657 22 315 649 DFFRX1 $T=55680 73660 0 180 $X=38260 $Y=67840
X256 658 13 12 659 22 315 592 DFFRX1 $T=56260 63220 1 180 $X=38840 $Y=62860
X257 660 13 12 661 22 315 662 DFFRX1 $T=69020 104980 0 180 $X=51600 $Y=99160
X258 596 13 12 663 22 315 590 DFFRX1 $T=69600 31900 1 180 $X=52180 $Y=31540
X259 664 13 12 665 22 315 666 DFFRX1 $T=71340 84100 1 180 $X=53920 $Y=83740
X260 667 13 12 668 22 315 669 DFFRX1 $T=72500 94540 1 180 $X=55080 $Y=94180
X261 670 13 12 671 22 24 35 DFFRX1 $T=62060 178060 1 0 $X=61460 $Y=172240
X262 672 13 12 31 22 24 673 DFFRX1 $T=80620 146740 1 180 $X=63200 $Y=146380
X263 674 13 12 675 22 24 676 DFFRX1 $T=83520 146740 0 180 $X=66100 $Y=140920
X264 677 13 12 678 22 315 679 DFFRX1 $T=88740 42340 1 180 $X=71320 $Y=41980
X265 42 13 12 41 22 24 39 DFFRX1 $T=96280 188500 0 180 $X=78860 $Y=182680
X266 680 13 12 40 22 24 681 DFFRX1 $T=100340 136300 1 180 $X=82920 $Y=135940
X267 629 13 12 628 22 24 682 DFFRX1 $T=102660 136300 0 180 $X=85240 $Y=130480
X268 683 13 12 684 22 24 44 DFFRX1 $T=85840 178060 0 0 $X=85240 $Y=177700
X269 685 13 12 686 22 24 687 DFFRX1 $T=103240 125860 0 180 $X=85820 $Y=120040
X270 688 13 12 689 22 315 595 DFFRX1 $T=106140 31900 0 180 $X=88720 $Y=26080
X271 690 13 12 691 22 315 602 DFFRX1 $T=106140 42340 0 180 $X=88720 $Y=36520
X272 692 13 12 693 22 315 677 DFFRX1 $T=106140 42340 1 180 $X=88720 $Y=41980
X273 694 13 12 695 22 315 696 DFFRX1 $T=106140 52780 1 180 $X=88720 $Y=52420
X274 697 13 12 698 22 315 699 DFFRX1 $T=89320 104980 1 0 $X=88720 $Y=99160
X275 700 13 12 701 22 24 702 DFFRX1 $T=106140 104980 1 180 $X=88720 $Y=104620
X276 703 13 12 704 22 315 601 DFFRX1 $T=125280 31900 0 180 $X=107860 $Y=26080
X277 705 13 12 48 22 24 706 DFFRX1 $T=125860 115420 1 180 $X=108440 $Y=115060
X278 707 13 12 30 22 24 50 DFFRX1 $T=125860 178060 1 180 $X=108440 $Y=177700
X279 708 13 12 709 22 24 56 DFFRX1 $T=113680 146740 1 0 $X=113080 $Y=140920
X280 710 13 12 711 22 24 52 DFFRX1 $T=131080 167620 1 180 $X=113660 $Y=167260
X281 712 13 12 713 22 320 714 DFFRX1 $T=125280 84100 0 0 $X=124680 $Y=83740
X282 715 13 12 716 22 24 63 DFFRX1 $T=125280 146740 0 0 $X=124680 $Y=146380
X283 717 13 12 718 22 320 719 DFFRX1 $T=143260 73660 1 180 $X=125840 $Y=73300
X284 720 13 12 721 22 320 722 DFFRX1 $T=143840 84100 0 180 $X=126420 $Y=78280
X285 723 13 12 724 22 320 725 DFFRX1 $T=144420 52780 0 180 $X=127000 $Y=46960
X286 726 13 12 727 22 320 728 DFFRX1 $T=144420 94540 0 180 $X=127000 $Y=88720
X287 729 13 12 64 22 320 730 DFFRX1 $T=148480 115420 0 180 $X=131060 $Y=109600
X288 731 13 12 732 22 24 67 DFFRX1 $T=141520 136300 0 0 $X=140920 $Y=135940
X289 733 13 12 734 22 320 606 DFFRX1 $T=164720 21460 1 180 $X=147300 $Y=21100
X290 735 13 12 736 22 320 703 DFFRX1 $T=165880 31900 0 180 $X=148460 $Y=26080
X291 737 13 12 738 22 320 739 DFFRX1 $T=173420 63220 1 180 $X=156000 $Y=62860
X292 740 13 12 741 22 320 742 DFFRX1 $T=157760 52780 1 0 $X=157160 $Y=46960
X293 68 13 12 743 22 24 69 DFFRX1 $T=176900 188500 0 180 $X=159480 $Y=182680
X294 77 13 12 72 22 320 744 DFFRX1 $T=178640 115420 1 180 $X=161220 $Y=115060
X295 745 13 12 746 22 320 747 DFFRX1 $T=180380 73660 0 180 $X=162960 $Y=67840
X296 748 13 12 749 22 320 750 DFFRX1 $T=180380 73660 1 180 $X=162960 $Y=73300
X297 751 13 12 632 22 320 752 DFFRX1 $T=187920 94540 0 180 $X=170500 $Y=88720
X298 753 13 12 754 22 320 755 DFFRX1 $T=187920 94540 1 180 $X=170500 $Y=94180
X299 756 13 12 757 22 320 758 DFFRX1 $T=194880 42340 0 180 $X=177460 $Y=36520
X300 759 13 12 760 22 320 761 DFFRX1 $T=195460 52780 0 180 $X=178040 $Y=46960
X301 762 13 12 763 22 24 80 DFFRX1 $T=179220 167620 1 0 $X=178620 $Y=161800
X302 764 13 12 765 22 85 87 DFFRX1 $T=198360 125860 0 0 $X=197760 $Y=125500
X303 766 13 12 767 22 24 88 DFFRX1 $T=198360 178060 0 0 $X=197760 $Y=177700
X304 768 13 12 769 22 85 733 DFFRX1 $T=215760 21460 1 180 $X=198340 $Y=21100
X305 770 13 12 771 22 85 772 DFFRX1 $T=220980 42340 0 180 $X=203560 $Y=36520
X306 773 13 12 774 22 85 83 DFFRX1 $T=222140 167620 0 180 $X=204720 $Y=161800
X307 79 13 12 93 22 85 775 DFFRX1 $T=222720 104980 0 180 $X=205300 $Y=99160
X308 776 13 12 777 22 85 611 DFFRX1 $T=226200 21460 0 180 $X=208780 $Y=15640
X309 778 13 12 779 22 85 780 DFFRX1 $T=229680 73660 1 180 $X=212260 $Y=73300
X310 781 13 12 782 22 85 783 DFFRX1 $T=230840 73660 0 180 $X=213420 $Y=67840
X311 784 13 12 785 22 85 786 DFFRX1 $T=232000 63220 0 180 $X=214580 $Y=57400
X312 787 13 12 788 22 85 789 DFFRX1 $T=238960 42340 0 180 $X=221540 $Y=36520
X313 790 13 12 791 22 85 792 DFFRX1 $T=241280 31900 1 180 $X=223860 $Y=31540
X314 793 13 12 794 22 85 795 DFFRX1 $T=242440 178060 1 180 $X=225020 $Y=177700
X315 796 13 12 797 22 85 798 DFFRX1 $T=243020 104980 0 180 $X=225600 $Y=99160
X316 98 13 12 799 22 85 38 DFFRX1 $T=244760 188500 0 180 $X=227340 $Y=182680
X317 615 13 12 800 22 85 776 DFFRX1 $T=245340 21460 0 180 $X=227920 $Y=15640
X318 801 13 12 33 22 85 802 DFFRX1 $T=247080 94540 0 180 $X=229660 $Y=88720
X319 803 13 12 804 22 85 805 DFFRX1 $T=259260 167620 1 180 $X=241840 $Y=167260
X320 806 13 12 807 22 85 100 DFFRX1 $T=262160 157180 0 180 $X=244740 $Y=151360
X321 808 13 12 809 22 85 810 DFFRX1 $T=263320 21460 1 180 $X=245900 $Y=21100
X322 811 13 12 812 22 85 101 DFFRX1 $T=266220 146740 1 180 $X=248800 $Y=146380
X323 813 13 12 814 22 85 102 DFFRX1 $T=266800 146740 0 180 $X=249380 $Y=140920
X324 815 13 12 816 22 85 103 DFFRX1 $T=269120 125860 1 180 $X=251700 $Y=125500
X325 817 13 12 818 22 85 107 DFFRX1 $T=262160 104980 1 0 $X=261560 $Y=99160
X326 819 13 12 820 22 85 821 DFFRX1 $T=263320 63220 0 0 $X=262720 $Y=62860
X327 822 13 12 823 22 85 824 DFFRX1 $T=265060 63220 1 0 $X=264460 $Y=57400
X328 825 13 12 826 22 85 827 DFFRX1 $T=284200 73660 0 180 $X=266780 $Y=67840
X329 828 13 12 829 22 85 111 DFFRX1 $T=269120 125860 0 0 $X=268520 $Y=125500
X330 830 13 12 831 22 118 832 DFFRX1 $T=305080 31900 1 180 $X=287660 $Y=31540
X331 833 13 12 834 22 118 835 DFFRX1 $T=305080 42340 0 180 $X=287660 $Y=36520
X332 836 13 12 837 22 118 838 DFFRX1 $T=305080 42340 1 180 $X=287660 $Y=41980
X333 839 13 12 840 22 118 841 DFFRX1 $T=305080 52780 0 180 $X=287660 $Y=46960
X334 842 13 12 843 22 118 844 DFFRX1 $T=305080 157180 0 180 $X=287660 $Y=151360
X335 845 13 12 846 22 118 847 DFFRX1 $T=305660 94540 1 180 $X=288240 $Y=94180
X336 848 13 12 849 22 118 850 DFFRX1 $T=307400 157180 1 180 $X=289980 $Y=156820
X337 851 13 12 852 22 118 853 DFFRX1 $T=307980 84100 1 180 $X=290560 $Y=83740
X338 854 13 12 855 22 118 856 DFFRX1 $T=307980 94540 0 180 $X=290560 $Y=88720
X339 857 13 12 858 22 118 859 DFFRX1 $T=319000 21460 1 180 $X=301580 $Y=21100
X340 860 13 12 861 22 118 862 DFFRX1 $T=324800 136300 1 180 $X=307380 $Y=135940
X341 863 13 12 864 22 118 865 DFFRX1 $T=326540 21460 0 180 $X=309120 $Y=15640
X342 124 13 12 108 22 118 866 DFFRX1 $T=326540 84100 1 180 $X=309120 $Y=83740
X343 867 13 12 868 22 118 869 DFFRX1 $T=327120 136300 0 180 $X=309700 $Y=130480
X344 870 13 12 871 22 118 872 DFFRX1 $T=338140 157180 1 180 $X=320720 $Y=156820
X345 873 13 12 874 22 118 875 DFFRX1 $T=339300 63220 1 180 $X=321880 $Y=62860
X346 876 13 12 877 22 118 878 DFFRX1 $T=339880 52780 1 180 $X=322460 $Y=52420
X347 879 13 12 880 22 118 881 DFFRX1 $T=339880 63220 0 180 $X=322460 $Y=57400
X348 882 13 12 883 22 118 884 DFFRX1 $T=339880 146740 1 180 $X=322460 $Y=146380
X349 885 13 12 886 22 118 887 DFFRX1 $T=341620 136300 1 180 $X=324200 $Y=135940
X350 888 13 12 889 22 118 890 DFFRX1 $T=346260 136300 0 180 $X=328840 $Y=130480
X351 621 13 12 891 22 118 614 DFFRX1 $T=348580 21460 1 180 $X=331160 $Y=21100
X352 892 13 12 893 22 118 894 DFFRX1 $T=354960 21460 0 180 $X=337540 $Y=15640
X353 895 13 12 896 22 118 897 DFFRX1 $T=358440 115420 1 180 $X=341020 $Y=115060
X354 898 13 12 899 22 118 900 DFFRX1 $T=358440 136300 1 180 $X=341020 $Y=135940
X355 901 13 12 902 22 118 903 DFFRX1 $T=362500 104980 1 180 $X=345080 $Y=104620
X356 134 13 12 135 22 118 904 DFFRX1 $T=352060 188500 1 0 $X=351460 $Y=182680
X357 905 13 12 906 22 118 907 DFFRX1 $T=369460 146740 1 180 $X=352040 $Y=146380
X358 908 13 12 909 22 118 910 DFFRX1 $T=372360 157180 0 180 $X=354940 $Y=151360
X359 138 13 12 137 22 118 911 DFFRX1 $T=375840 73660 0 180 $X=358420 $Y=67840
X360 140 13 12 143 22 118 912 DFFRX1 $T=378160 188500 1 0 $X=377560 $Y=182680
X361 913 13 12 914 22 474 915 DFFRX1 $T=398460 73660 0 180 $X=381040 $Y=67840
X362 916 13 12 917 22 118 918 DFFRX1 $T=383380 157180 1 0 $X=382780 $Y=151360
X363 919 13 12 920 22 474 921 DFFRX1 $T=404260 63220 1 180 $X=386840 $Y=62860
X364 922 13 12 923 22 474 924 DFFRX1 $T=406000 73660 1 180 $X=388580 $Y=73300
X365 925 13 12 926 22 474 927 DFFRX1 $T=408320 42340 1 180 $X=390900 $Y=41980
X366 152 13 12 151 22 474 928 DFFRX1 $T=413540 104980 0 180 $X=396120 $Y=99160
X367 929 13 12 930 22 474 931 DFFRX1 $T=414700 104980 1 180 $X=397280 $Y=104620
X368 932 13 12 933 22 474 934 DFFRX1 $T=417020 42340 0 180 $X=399600 $Y=36520
X369 935 13 12 936 22 474 937 DFFRX1 $T=419340 31900 0 180 $X=401920 $Y=26080
X370 146 13 12 150 22 141 938 DFFRX1 $T=404260 188500 1 0 $X=403660 $Y=182680
X371 939 13 12 940 22 141 941 DFFRX1 $T=405420 167620 1 0 $X=404820 $Y=161800
X372 942 13 12 943 22 474 944 DFFRX1 $T=432680 125860 1 180 $X=415260 $Y=125500
X373 945 13 12 946 22 141 947 DFFRX1 $T=432680 146740 1 180 $X=415260 $Y=146380
X374 948 13 12 949 22 474 950 DFFRX1 $T=433840 115420 1 180 $X=416420 $Y=115060
X375 159 13 12 154 22 141 951 DFFRX1 $T=439060 188500 0 180 $X=421640 $Y=182680
X376 952 13 12 953 22 474 618 DFFRX1 $T=439640 21460 0 180 $X=422220 $Y=15640
X377 954 13 12 955 22 474 956 DFFRX1 $T=439640 63220 0 180 $X=422220 $Y=57400
X378 957 13 12 958 22 474 959 DFFRX1 $T=440220 52780 1 180 $X=422800 $Y=52420
X379 960 13 12 961 22 474 962 DFFRX1 $T=441380 42340 0 180 $X=423960 $Y=36520
X380 963 13 12 964 22 474 965 DFFRX1 $T=441960 63220 1 180 $X=424540 $Y=62860
X381 966 13 12 967 22 474 968 DFFRX1 $T=442540 52780 0 180 $X=425120 $Y=46960
X382 969 13 12 970 22 474 971 DFFRX1 $T=443700 73660 1 180 $X=426280 $Y=73300
X383 972 13 12 973 22 474 974 DFFRX1 $T=443700 84100 1 180 $X=426280 $Y=83740
X384 975 13 12 976 22 474 977 DFFRX1 $T=444280 84100 0 180 $X=426860 $Y=78280
X385 167 13 12 162 22 474 978 DFFRX1 $T=452400 104980 1 180 $X=434980 $Y=104620
X386 168 13 12 165 22 141 979 DFFRX1 $T=458200 157180 0 180 $X=440780 $Y=151360
X387 980 13 12 981 22 474 624 DFFRX1 $T=458780 21460 0 180 $X=441360 $Y=15640
X388 982 13 12 983 22 141 984 DFFRX1 $T=464000 115420 1 180 $X=446580 $Y=115060
X389 985 13 12 986 22 141 987 DFFRX1 $T=464580 136300 1 180 $X=447160 $Y=135940
X390 988 13 12 989 22 141 990 DFFRX1 $T=464580 146740 0 180 $X=447160 $Y=140920
X391 991 13 12 992 22 141 952 DFFRX1 $T=484880 21460 0 180 $X=467460 $Y=15640
X392 993 13 12 994 22 141 995 DFFRX1 $T=484880 31900 0 180 $X=467460 $Y=26080
X393 996 13 12 997 22 141 998 DFFRX1 $T=484880 42340 0 180 $X=467460 $Y=36520
X394 999 13 12 1000 22 141 1001 DFFRX1 $T=484880 52780 0 180 $X=467460 $Y=46960
X395 1002 13 12 1003 22 141 1004 DFFRX1 $T=484880 52780 1 180 $X=467460 $Y=52420
X396 1005 13 12 1006 22 141 1007 DFFRX1 $T=484880 63220 0 180 $X=467460 $Y=57400
X397 1008 13 12 1009 22 141 1010 DFFRX1 $T=484880 73660 0 180 $X=467460 $Y=67840
X398 1011 13 12 1012 22 141 1013 DFFRX1 $T=484880 84100 0 180 $X=467460 $Y=78280
X399 1014 13 12 1015 22 141 1016 DFFRX1 $T=484880 94540 1 180 $X=467460 $Y=94180
X400 1017 13 12 1018 22 141 1019 DFFRX1 $T=468640 146740 1 0 $X=468040 $Y=140920
X401 1020 13 12 1021 22 141 1022 DFFRX1 $T=473280 104980 0 0 $X=472680 $Y=104620
X402 1023 13 12 1024 22 141 1025 DFFRX1 $T=483140 84100 0 0 $X=482540 $Y=83740
X403 1026 13 12 184 22 141 1027 DFFRX1 $T=500540 167620 1 180 $X=483120 $Y=167260
X404 180 13 12 185 22 141 1028 DFFRX1 $T=500540 178060 1 180 $X=483120 $Y=177700
X405 1029 13 12 1030 22 141 1031 DFFRX1 $T=504600 136300 1 180 $X=487180 $Y=135940
X406 1032 13 12 1033 22 141 1034 DFFRX1 $T=505760 125860 1 180 $X=488340 $Y=125500
X407 1035 13 12 1036 22 141 1037 DFFRX1 $T=506340 115420 1 180 $X=488920 $Y=115060
X408 181 13 12 1038 22 141 1039 DFFRX1 $T=506340 167620 0 180 $X=488920 $Y=161800
X409 186 13 12 183 22 141 1040 DFFRX1 $T=509240 104980 0 180 $X=491820 $Y=99160
X410 1041 13 12 1042 22 141 1043 DFFRX1 $T=509820 52780 0 180 $X=492400 $Y=46960
X411 1044 13 12 1045 22 141 1046 DFFRX1 $T=509820 63220 0 180 $X=492400 $Y=57400
X412 1047 13 12 1048 22 141 1049 DFFRX1 $T=509820 94540 1 180 $X=492400 $Y=94180
X413 1050 13 12 1051 22 141 1052 DFFRX1 $T=512720 73660 1 180 $X=495300 $Y=73300
X414 1053 13 12 1054 22 141 1055 DFFRX1 $T=513300 63220 1 180 $X=495880 $Y=62860
X415 193 13 12 189 22 141 1056 DFFRX1 $T=513880 157180 0 180 $X=496460 $Y=151360
X416 1057 13 12 1058 22 141 1059 DFFRX1 $T=516780 42340 0 180 $X=499360 $Y=36520
X417 1060 13 12 1061 22 141 1062 DFFRX1 $T=516780 84100 1 180 $X=499360 $Y=83740
X418 190 13 12 1063 22 141 1064 DFFRX1 $T=510980 157180 0 0 $X=510380 $Y=156820
X419 1065 13 12 1066 22 141 1067 DFFRX1 $T=534180 115420 1 180 $X=516760 $Y=115060
X420 1068 13 12 1069 22 141 1070 DFFRX1 $T=535920 104980 1 180 $X=518500 $Y=104620
X421 1071 13 12 1072 22 141 625 DFFRX1 $T=537080 21460 1 180 $X=519660 $Y=21100
X422 1073 13 12 1074 22 141 1075 DFFRX1 $T=537660 31900 1 180 $X=520240 $Y=31540
X423 1076 13 12 1077 22 141 1078 DFFRX1 $T=537660 63220 1 180 $X=520240 $Y=62860
X424 1079 13 12 1080 22 141 1081 DFFRX1 $T=537660 73660 1 180 $X=520240 $Y=73300
X425 1082 13 12 1083 22 141 1084 DFFRX1 $T=537660 84100 1 180 $X=520240 $Y=83740
X426 1085 13 12 1086 22 141 1087 DFFRX1 $T=537660 94540 0 180 $X=520240 $Y=88720
X427 1088 13 12 1089 22 141 1090 DFFRX1 $T=538240 42340 1 180 $X=520820 $Y=41980
X428 1091 13 12 1092 22 141 1093 DFFRX1 $T=541720 63220 0 180 $X=524300 $Y=57400
X429 1094 13 12 1095 22 24 639 227 640 SDFFRXL $T=71920 115420 1 180 $X=50440 $Y=115060
X430 1096 13 12 1097 22 24 644 1098 643 SDFFRXL $T=72500 125860 1 180 $X=51020 $Y=125500
X431 1099 13 12 1100 22 315 657 1101 656 SDFFRXL $T=73660 73660 1 180 $X=52180 $Y=73300
X432 1102 13 12 1103 22 24 1095 1104 1094 SDFFRXL $T=81780 115420 0 180 $X=60300 $Y=109600
X433 1105 13 12 1106 22 315 658 239 659 SDFFRXL $T=83520 63220 1 180 $X=62040 $Y=62860
X434 1107 13 12 1108 22 315 664 241 665 SDFFRXL $T=83520 84100 0 180 $X=62040 $Y=78280
X435 1109 13 12 1110 22 315 668 1111 667 SDFFRXL $T=84680 94540 0 180 $X=63200 $Y=88720
X436 1112 13 12 1113 22 315 1106 1114 1105 SDFFRXL $T=106140 63220 1 180 $X=84660 $Y=62860
X437 1115 13 12 1116 22 315 1099 255 1100 SDFFRXL $T=106140 73660 0 180 $X=84660 $Y=67840
X438 1117 13 12 1118 22 315 1108 1119 1107 SDFFRXL $T=106140 84100 0 180 $X=84660 $Y=78280
X439 1120 13 12 1121 22 315 698 1122 697 SDFFRXL $T=106140 94540 1 180 $X=84660 $Y=94180
X440 1123 13 12 1124 22 24 686 1125 685 SDFFRXL $T=106140 115420 0 180 $X=84660 $Y=109600
X441 1126 13 12 1127 22 24 257 45 46 SDFFRXL $T=85260 167620 0 0 $X=84660 $Y=167260
X442 1128 13 12 1129 22 320 689 1130 688 SDFFRXL $T=131080 31900 1 180 $X=109600 $Y=31540
X443 1131 13 12 1132 22 24 55 59 266 SDFFRXL $T=113100 167620 1 0 $X=112500 $Y=161800
X444 1133 13 12 1134 22 320 1116 1135 1115 SDFFRXL $T=141520 63220 1 180 $X=120040 $Y=62860
X445 1136 13 12 1137 22 320 1124 1138 1123 SDFFRXL $T=145580 104980 0 180 $X=124100 $Y=99160
X446 1139 13 12 1140 22 320 1112 272 1113 SDFFRXL $T=147900 63220 0 180 $X=126420 $Y=57400
X447 1141 13 12 1142 22 320 701 1143 700 SDFFRXL $T=147900 94540 1 180 $X=126420 $Y=94180
X448 1144 13 12 1145 22 320 274 627 273 SDFFRXL $T=150800 115420 1 180 $X=129320 $Y=115060
X449 1146 13 12 1147 22 320 277 48 276 SDFFRXL $T=151960 31900 1 180 $X=130480 $Y=31540
X450 1148 13 12 1149 22 320 1140 1150 1139 SDFFRXL $T=180960 63220 0 180 $X=159480 $Y=57400
X451 1151 13 12 1152 22 320 727 1153 726 SDFFRXL $T=182700 84100 1 180 $X=161220 $Y=83740
X452 1154 13 12 1155 22 320 1147 1156 1146 SDFFRXL $T=184440 31900 1 180 $X=162960 $Y=31540
X453 1157 13 12 1158 22 320 319 1137 318 SDFFRXL $T=189660 104980 0 180 $X=168180 $Y=99160
X454 1159 13 12 1160 22 320 740 317 741 SDFFRXL $T=190820 52780 1 180 $X=169340 $Y=52420
X455 1161 13 12 1162 22 24 76 74 321 SDFFRXL $T=190820 167620 1 180 $X=169340 $Y=167260
X456 1163 13 12 1164 22 85 343 330 84 SDFFRXL $T=219240 167620 1 180 $X=197760 $Y=167260
X457 1165 13 12 1166 22 85 350 94 86 SDFFRXL $T=199520 178060 1 0 $X=198920 $Y=172240
X458 1167 13 12 1168 22 85 1158 1169 1157 SDFFRXL $T=226200 84100 1 180 $X=204720 $Y=83740
X459 1170 13 12 1171 22 85 754 1172 753 SDFFRXL $T=226200 94540 0 180 $X=204720 $Y=88720
X460 1173 13 12 1174 22 85 759 346 760 SDFFRXL $T=231420 52780 0 180 $X=209940 $Y=46960
X461 1175 13 12 1176 22 85 1160 1177 1159 SDFFRXL $T=233740 52780 1 180 $X=212260 $Y=52420
X462 97 13 12 96 22 85 368 1178 367 SDFFRXL $T=241280 178060 0 180 $X=219800 $Y=172240
X463 1179 13 12 1180 22 85 363 356 364 SDFFRXL $T=241860 167620 1 180 $X=220380 $Y=167260
X464 1181 13 12 1182 22 85 375 72 376 SDFFRXL $T=247080 31900 0 180 $X=225600 $Y=26080
X465 635 13 12 634 22 85 1171 1183 1170 SDFFRXL $T=251140 84100 1 180 $X=229660 $Y=83740
X466 1184 13 12 1185 22 85 1168 1186 1167 SDFFRXL $T=270280 84100 0 180 $X=248800 $Y=78280
X467 1187 13 12 1188 22 85 402 631 401 SDFFRXL $T=278980 73660 1 180 $X=257500 $Y=73300
X468 865 13 12 1189 22 85 93 394 79 SDFFRXL $T=283040 21460 0 180 $X=261560 $Y=15640
X469 1190 13 12 1191 22 85 406 809 405 SDFFRXL $T=284200 21460 1 180 $X=262720 $Y=21100
X470 1192 13 12 1193 22 85 819 408 820 SDFFRXL $T=284200 52780 0 180 $X=262720 $Y=46960
X471 1194 13 12 1195 22 85 823 1196 822 SDFFRXL $T=284200 52780 1 180 $X=262720 $Y=52420
X472 116 13 12 115 22 118 420 1197 421 SDFFRXL $T=309140 146740 1 180 $X=287660 $Y=146380
X473 1198 13 12 1199 22 118 425 1200 424 SDFFRXL $T=319580 104980 0 180 $X=298100 $Y=99160
X474 1201 13 12 1202 22 118 431 1203 430 SDFFRXL $T=328280 115420 1 180 $X=306800 $Y=115060
X475 1204 13 12 1205 22 118 1193 1206 1192 SDFFRXL $T=333500 52780 0 180 $X=312020 $Y=46960
X476 1207 13 12 1208 22 118 439 852 438 SDFFRXL $T=335240 73660 1 180 $X=313760 $Y=73300
X477 1209 13 12 1210 22 118 440 420 441 SDFFRXL $T=338140 146740 0 180 $X=316660 $Y=140920
X478 1211 13 12 1212 22 118 858 1213 857 SDFFRXL $T=341620 31900 0 180 $X=320140 $Y=26080
X479 1214 13 12 1215 22 118 436 837 437 SDFFRXL $T=341620 42340 0 180 $X=320140 $Y=36520
X480 1216 13 12 1217 22 118 442 831 443 SDFFRXL $T=342200 31900 1 180 $X=320720 $Y=31540
X481 1218 13 12 1219 22 118 834 445 833 SDFFRXL $T=342780 42340 1 180 $X=321300 $Y=41980
X482 1220 13 12 1221 22 118 447 1185 446 SDFFRXL $T=343940 84100 0 180 $X=322460 $Y=78280
X483 1222 13 12 1223 22 474 466 1212 467 SDFFRXL $T=375840 21460 0 180 $X=354360 $Y=15640
X484 937 13 12 1224 22 474 463 893 462 SDFFRXL $T=375840 31900 0 180 $X=354360 $Y=26080
X485 1225 13 12 1226 22 474 464 1217 465 SDFFRXL $T=375840 31900 1 180 $X=354360 $Y=31540
X486 1227 13 12 1228 22 474 468 1219 469 SDFFRXL $T=375840 52780 0 180 $X=354360 $Y=46960
X487 1229 13 12 1230 22 118 460 1215 461 SDFFRXL $T=375840 52780 1 180 $X=354360 $Y=52420
X488 142 13 12 144 22 118 472 1231 473 SDFFRXL $T=399040 178060 0 180 $X=377560 $Y=172240
X489 1232 13 12 1233 22 474 476 616 475 SDFFRXL $T=399620 84100 0 180 $X=378140 $Y=78280
X490 1234 13 12 1235 22 474 1221 1236 1220 SDFFRXL $T=400200 84100 1 180 $X=378720 $Y=83740
X491 1237 13 12 1238 22 474 477 633 478 SDFFRXL $T=400780 94540 0 180 $X=379300 $Y=88720
X492 149 13 12 148 22 141 497 1231 498 SDFFRXL $T=406000 178060 1 180 $X=384520 $Y=177700
X493 1239 13 12 1240 22 474 1238 1241 1237 SDFFRXL $T=417600 94540 1 180 $X=396120 $Y=94180
X494 1242 13 12 1243 22 474 520 1233 519 SDFFRXL $T=434420 104980 0 180 $X=412940 $Y=99160
X495 1244 13 12 1245 22 474 525 1235 526 SDFFRXL $T=436160 94540 0 180 $X=414680 $Y=88720
X496 1246 13 12 1247 22 474 137 1248 138 SDFFRXL $T=436740 31900 1 180 $X=415260 $Y=31540
X497 1249 13 12 1250 22 474 1243 1251 1242 SDFFRXL $T=462840 115420 0 180 $X=441360 $Y=109600
X498 1252 13 12 1253 22 141 151 1254 152 SDFFRXL $T=488940 31900 1 180 $X=467460 $Y=31540
X499 1255 13 12 1256 22 141 556 1240 555 SDFFRXL $T=488940 104980 0 180 $X=467460 $Y=99160
X500 1257 13 12 1258 22 141 1256 1259 1255 SDFFRXL $T=506920 115420 0 180 $X=485440 $Y=109600
X501 1075 13 12 1260 22 141 568 1253 567 SDFFRXL $T=513300 31900 1 180 $X=491820 $Y=31540
X502 1261 13 12 1262 22 141 571 994 572 SDFFRXL $T=516200 21460 1 180 $X=494720 $Y=21100
X503 1263 13 12 1264 22 141 1258 1265 1257 SDFFRXL $T=517940 146740 1 180 $X=496460 $Y=146380
X504 1266 13 12 1267 22 141 580 1030 579 SDFFRXL $T=530120 146740 0 180 $X=508640 $Y=140920
X505 1268 13 12 1269 22 141 584 1033 583 SDFFRXL $T=531280 125860 0 180 $X=509800 $Y=120040
X506 1270 13 12 1271 22 141 186 1272 183 SDFFRXL $T=541140 42340 0 180 $X=519660 $Y=36520
X507 711 670 13 12 1273 795 XNOR3X1 $T=78880 178060 1 0 $X=78280 $Y=172240
X508 1127 683 13 12 1274 805 XNOR3X1 $T=84100 167620 1 0 $X=83500 $Y=161800
X509 599 677 13 12 40 696 XNOR3X1 $T=88740 52780 1 0 $X=88140 $Y=46960
X510 1132 708 13 12 1275 844 XNOR3X1 $T=115420 157180 1 0 $X=114820 $Y=151360
X511 732 715 13 12 1276 884 XNOR3X1 $T=132820 146740 1 0 $X=132220 $Y=140920
X512 736 733 13 12 729 772 XNOR3X1 $T=162400 42340 0 0 $X=161800 $Y=41980
X513 732 53 13 12 1277 850 XNOR3X1 $T=167040 146740 0 0 $X=166440 $Y=146380
X514 607 1161 13 12 1278 887 XNOR3X1 $T=172260 136300 0 0 $X=171660 $Y=135940
X515 743 49 13 12 1279 82 XNOR3X1 $T=178640 188500 1 0 $X=178040 $Y=182680
X516 1164 766 13 12 1280 869 XNOR3X1 $T=198360 136300 1 0 $X=197760 $Y=130480
X517 765 1165 13 12 1281 847 XNOR3X1 $T=204740 115420 0 0 $X=204140 $Y=115060
X518 763 773 13 12 1282 872 XNOR3X1 $T=207640 157180 0 0 $X=207040 $Y=156820
X519 774 1162 13 12 1283 862 XNOR3X1 $T=227360 146740 0 0 $X=226760 $Y=146380
X520 807 1161 13 12 1284 918 XNOR3X1 $T=251720 157180 1 180 $X=233720 $Y=156820
X521 804 1179 13 12 1285 109 XNOR3X1 $T=263320 167620 0 0 $X=262720 $Y=167260
X522 797 817 13 12 1286 856 XNOR3X1 $T=263900 94540 1 0 $X=263300 $Y=88720
X523 815 1162 13 12 1287 900 XNOR3X1 $T=267380 125860 1 0 $X=266780 $Y=120040
X524 811 1162 13 12 1288 910 XNOR3X1 $T=268540 146740 1 0 $X=267940 $Y=140920
X525 1189 1190 13 12 801 894 XNOR3X1 $T=288260 21460 1 0 $X=287660 $Y=15640
X526 829 815 13 12 1289 903 XNOR3X1 $T=288260 125860 1 0 $X=287660 $Y=120040
X527 96 793 13 12 1290 114 XNOR3X1 $T=288260 178060 0 0 $X=287660 $Y=177700
X528 812 813 13 12 1291 890 XNOR3X1 $T=291740 136300 1 0 $X=291140 $Y=130480
X529 849 115 13 12 1292 904 XNOR3X1 $T=316100 178060 1 0 $X=315500 $Y=172240
X530 849 842 13 12 1293 912 XNOR3X1 $T=317260 167620 0 0 $X=316660 $Y=167260
X531 846 1201 13 12 1294 931 XNOR3X1 $T=327700 104980 0 0 $X=327100 $Y=104620
X532 871 115 13 12 1295 130 XNOR3X1 $T=330020 167620 1 0 $X=329420 $Y=161800
X533 883 1210 13 12 1296 136 XNOR3X1 $T=342200 178060 1 0 $X=341600 $Y=172240
X534 886 1210 13 12 1297 938 XNOR3X1 $T=344520 167620 0 0 $X=343920 $Y=167260
X535 1199 854 13 12 1298 944 XNOR3X1 $T=345100 94540 0 0 $X=344500 $Y=94180
X536 861 867 13 12 1299 941 XNOR3X1 $T=348000 136300 1 0 $X=347400 $Y=130480
X537 899 888 13 12 1300 1019 XNOR3X1 $T=358440 136300 0 0 $X=357840 $Y=135940
X538 896 901 13 12 1301 984 XNOR3X1 $T=378160 104980 1 0 $X=377560 $Y=99160
X539 916 1210 13 12 1302 145 XNOR3X1 $T=379320 167620 1 0 $X=378720 $Y=161800
X540 864 621 13 12 124 619 XNOR3X1 $T=379900 21460 0 0 $X=379300 $Y=21100
X541 861 1210 13 12 1303 947 XNOR3X1 $T=390340 146740 1 0 $X=389740 $Y=140920
X542 908 1210 13 12 1304 951 XNOR3X1 $T=390340 157180 0 0 $X=389740 $Y=156820
X543 898 1210 13 12 1305 979 XNOR3X1 $T=395560 146740 0 0 $X=394960 $Y=146380
X544 940 149 13 12 1306 155 XNOR3X1 $T=412380 178060 0 0 $X=411780 $Y=177700
X545 946 144 13 12 1307 161 XNOR3X1 $T=433840 157180 0 0 $X=433240 $Y=156820
X546 946 929 13 12 1308 163 XNOR3X1 $T=435000 146740 0 0 $X=434400 $Y=146380
X547 949 942 13 12 1309 1064 XNOR3X1 $T=437900 136300 1 0 $X=437300 $Y=130480
X548 986 982 13 12 1310 1039 XNOR3X1 $T=468060 136300 0 0 $X=467460 $Y=135940
X549 1018 988 13 12 1311 1027 XNOR3X1 $T=468060 167620 1 0 $X=467460 $Y=161800
X550 992 980 13 12 162 626 XNOR3X1 $T=484880 21460 1 0 $X=484280 $Y=15640
X551 640 13 12 653 23 1098 639 228 OAI221XL $T=55680 125860 1 0 $X=55080 $Y=120040
X552 659 13 12 31 672 1101 658 238 OAI221XL $T=70760 63220 0 180 $X=64360 $Y=57400
X553 665 13 12 31 672 1111 664 240 OAI221XL $T=71340 84100 0 0 $X=70740 $Y=83740
X554 1106 13 12 40 680 255 1105 1114 OAI221XL $T=90480 73660 1 180 $X=84080 $Y=73300
X555 1100 13 12 40 680 1119 1099 256 OAI221XL $T=95120 73660 0 0 $X=94520 $Y=73300
X556 691 13 12 48 705 1130 703 268 OAI221XL $T=124700 42340 0 180 $X=118300 $Y=36520
X557 1112 13 12 48 705 1135 1113 271 OAI221XL $T=121220 63220 1 0 $X=120620 $Y=57400
X558 741 13 12 729 64 1150 740 316 OAI221XL $T=164720 52780 1 180 $X=158320 $Y=52420
X559 759 13 12 72 77 1177 760 347 OAI221XL $T=212860 52780 1 180 $X=206460 $Y=52420
X560 820 13 12 93 79 1196 819 407 OAI221XL $T=264480 42340 0 0 $X=263880 $Y=41980
X561 1312 13 12 1313 116 1314 848 1315 OAI221XL $T=310300 178060 1 0 $X=309700 $Y=172240
X562 837 13 12 33 801 1206 836 436 OAI221XL $T=320160 42340 1 180 $X=313760 $Y=41980
X563 858 13 12 801 33 442 857 1213 OAI221XL $T=319580 21460 0 0 $X=318980 $Y=21100
X564 128 13 12 116 452 131 132 457 OAI221XL $T=343940 188500 1 0 $X=343340 $Y=182680
X565 892 13 12 108 124 466 893 463 OAI221XL $T=357860 21460 0 0 $X=357260 $Y=21100
X566 1219 13 12 108 124 460 1218 468 OAI221XL $T=363080 42340 0 0 $X=362480 $Y=41980
X567 860 13 12 1209 1316 1317 1318 1319 OAI221XL $T=381640 115420 0 0 $X=381040 $Y=115060
X568 945 13 12 142 1320 1321 1322 1323 OAI221XL $T=435000 178060 0 0 $X=434400 $Y=177700
X569 1253 13 12 162 167 571 1252 568 OAI221XL $T=494740 31900 1 0 $X=494140 $Y=26080
X570 1324 642 13 12 646 223 OR3X1 $T=45820 115420 1 0 $X=45220 $Y=109600
X571 1325 641 13 12 645 1326 OR3X1 $T=53360 104980 0 0 $X=52760 $Y=104620
X572 1327 660 13 12 1094 234 OR3X1 $T=60900 104980 0 0 $X=60300 $Y=104620
X573 1328 692 13 12 694 1329 OR3X1 $T=99760 63220 1 0 $X=99160 $Y=57400
X574 1330 693 13 12 695 1331 OR3X1 $T=111360 52780 1 0 $X=110760 $Y=46960
X575 1332 700 13 12 1123 264 OR3X1 $T=116580 104980 0 0 $X=115980 $Y=104620
X576 1333 701 13 12 1121 1334 OR3X1 $T=121800 94540 0 0 $X=121200 $Y=94180
X577 1335 1129 13 12 724 299 OR3X1 $T=142100 42340 0 0 $X=141500 $Y=41980
X578 1336 1128 13 12 723 1337 OR3X1 $T=151380 52780 0 180 $X=146140 $Y=46960
X579 1338 64 13 12 721 1339 OR3X1 $T=150220 84100 0 0 $X=149620 $Y=83740
X580 1340 745 13 12 748 1341 OR3X1 $T=180960 73660 0 0 $X=180360 $Y=73300
X581 1342 785 13 12 782 369 OR3X1 $T=236640 63220 1 180 $X=231400 $Y=62860
X582 369 631 13 12 779 1343 OR3X1 $T=232000 73660 0 0 $X=231400 $Y=73300
X583 1344 784 13 12 781 1345 OR3X1 $T=238960 63220 0 0 $X=238360 $Y=62860
X584 1346 1173 13 12 1175 397 OR3X1 $T=249980 42340 0 0 $X=249380 $Y=41980
X585 418 33 13 12 826 1347 OR3X1 $T=293480 73660 1 0 $X=292880 $Y=67840
X586 1348 1195 13 12 840 418 OR3X1 $T=298700 52780 1 180 $X=293460 $Y=52420
X587 1349 1194 13 12 839 1350 OR3X1 $T=299280 63220 0 180 $X=294040 $Y=57400
X588 1351 880 13 12 874 458 OR3X1 $T=339300 63220 0 0 $X=338700 $Y=62860
X589 1352 1205 13 12 877 1351 OR3X1 $T=342200 52780 0 0 $X=341600 $Y=52420
X590 1353 1204 13 12 876 1354 OR3X1 $T=353220 52780 1 180 $X=347980 $Y=52420
X591 1354 879 13 12 873 1355 OR3X1 $T=353220 63220 1 180 $X=347980 $Y=62860
X592 458 616 13 12 1208 1356 OR3X1 $T=361340 73660 0 0 $X=360740 $Y=73300
X593 1357 1227 13 12 1229 1358 OR3X1 $T=397880 52780 0 0 $X=397280 $Y=52420
X594 1359 919 13 12 913 1360 OR3X1 $T=403100 73660 1 0 $X=402500 $Y=67840
X595 506 491 13 12 1361 1362 OR3X1 $T=403100 115420 0 0 $X=402500 $Y=115060
X596 1358 925 13 12 932 1359 OR3X1 $T=410640 52780 0 0 $X=410040 $Y=52420
X597 1363 957 13 12 954 1364 OR3X1 $T=443700 63220 0 0 $X=443100 $Y=62860
X598 1365 960 13 12 966 1363 OR3X1 $T=450660 42340 1 180 $X=445420 $Y=41980
X599 1364 963 13 12 969 1366 OR3X1 $T=457040 73660 0 180 $X=451800 $Y=67840
X600 560 542 13 12 1367 1368 OR3X1 $T=468060 167620 0 0 $X=467460 $Y=167260
X601 1369 1020 13 12 1249 1370 OR3X1 $T=475020 115420 0 180 $X=469780 $Y=109600
X602 1371 996 13 12 999 1372 OR3X1 $T=477340 42340 1 180 $X=472100 $Y=41980
X603 1372 1002 13 12 1005 1373 OR3X1 $T=472700 63220 0 0 $X=472100 $Y=62860
X604 1374 1023 13 12 1014 1369 OR3X1 $T=480820 94540 0 180 $X=475580 $Y=88720
X605 1375 1009 13 12 1012 1376 OR3X1 $T=483720 73660 1 180 $X=478480 $Y=73300
X606 1377 997 13 12 1000 1378 OR3X1 $T=484880 52780 1 0 $X=484280 $Y=46960
X607 1378 1003 13 12 1006 1375 OR3X1 $T=489520 63220 0 180 $X=484280 $Y=57400
X608 1373 1008 13 12 1011 1374 OR3X1 $T=489520 73660 1 180 $X=484280 $Y=73300
X609 1376 1024 13 12 1015 557 OR3X1 $T=489520 94540 1 180 $X=484280 $Y=94180
X610 576 1033 13 12 1036 1379 OR3X1 $T=502280 125860 0 180 $X=497040 $Y=120040
X611 1380 1060 13 12 1047 1381 OR3X1 $T=510400 104980 0 0 $X=509800 $Y=104620
X612 1382 1053 13 12 1050 1380 OR3X1 $T=518520 73660 1 180 $X=513280 $Y=73300
X613 707 13 12 1383 53 282 1384 OAI211XL $T=133980 178060 1 0 $X=133380 $Y=172240
X614 815 13 12 1385 1162 389 1386 OAI211XL $T=252880 115420 0 0 $X=252280 $Y=115060
X615 898 13 12 1387 1210 481 500 OAI211XL $T=393820 136300 0 0 $X=393220 $Y=135940
X616 672 13 12 230 236 1388 237 31 OAI32XL $T=69020 52780 0 180 $X=63200 $Y=46960
X617 660 13 12 31 1327 1104 1389 672 OAI32XL $T=65540 104980 0 0 $X=64940 $Y=104620
X618 1109 13 12 40 253 1122 1390 680 OAI32XL $T=89900 94540 0 180 $X=84080 $Y=88720
X619 1391 13 12 310 314 363 1392 801 OAI32XL $T=166460 167620 0 180 $X=160640 $Y=161800
X620 1393 13 12 378 366 1203 1394 33 OAI32XL $T=240120 125860 0 0 $X=239520 $Y=125500
X621 1250 13 12 1021 1395 1259 1370 167 OAI32XL $T=475020 115420 1 0 $X=474420 $Y=109600
X622 1324 13 12 653 1396 OR2X1 $T=44660 115420 0 180 $X=40580 $Y=109600
X623 1325 13 12 23 1397 OR2X1 $T=53360 104980 1 180 $X=49280 $Y=104620
X624 663 13 12 648 229 OR2X1 $T=62060 42340 0 180 $X=57980 $Y=36520
X625 1398 13 12 661 1389 OR2X1 $T=74240 104980 1 180 $X=70160 $Y=104620
X626 1388 13 12 1399 679 OR2X1 $T=71340 52780 1 0 $X=70740 $Y=46960
X627 1400 13 12 1096 1401 OR2X1 $T=77720 125860 1 180 $X=73640 $Y=125500
X628 1402 13 12 1110 1390 OR2X1 $T=80040 84100 0 0 $X=79440 $Y=83740
X629 1403 13 12 1103 1404 OR2X1 $T=81780 115420 1 0 $X=81180 $Y=109600
X630 678 13 12 599 244 OR2X1 $T=83520 52780 0 0 $X=82920 $Y=52420
X631 1390 13 12 698 246 OR2X1 $T=85840 104980 1 0 $X=85240 $Y=99160
X632 1405 13 12 1120 1332 OR2X1 $T=110780 94540 0 0 $X=110180 $Y=94180
X633 1330 13 12 48 1406 OR2X1 $T=120060 52780 0 180 $X=115980 $Y=46960
X634 1328 13 12 705 1407 OR2X1 $T=116580 63220 1 0 $X=115980 $Y=57400
X635 259 13 12 705 1408 OR2X1 $T=117160 73660 1 0 $X=116560 $Y=67840
X636 49 13 12 41 1409 OR2X1 $T=118320 188500 1 0 $X=117720 $Y=182680
X637 263 13 12 48 1410 OR2X1 $T=121800 73660 1 0 $X=121200 $Y=67840
X638 1334 13 12 48 1411 OR2X1 $T=125860 104980 1 180 $X=121780 $Y=104620
X639 1412 13 12 53 282 OR2X1 $T=138620 178060 1 180 $X=134540 $Y=177700
X640 1335 13 12 64 1413 OR2X1 $T=136300 42340 0 0 $X=135700 $Y=41980
X641 1127 13 12 1132 1414 OR2X1 $T=136300 157180 1 0 $X=135700 $Y=151360
X642 1412 13 12 49 295 OR2X1 $T=138620 188500 1 0 $X=138020 $Y=182680
X643 711 13 12 30 1415 OR2X1 $T=141520 167620 0 0 $X=140920 $Y=167260
X644 53 13 12 732 1416 OR2X1 $T=144420 146740 0 0 $X=143820 $Y=146380
X645 1417 13 12 720 1418 OR2X1 $T=145000 84100 0 0 $X=144400 $Y=83740
X646 1419 13 12 1420 1178 OR2X1 $T=149640 167620 1 0 $X=149040 $Y=161800
X647 1418 13 12 729 301 OR2X1 $T=151380 94540 0 0 $X=150780 $Y=94180
X648 294 13 12 729 1421 OR2X1 $T=151960 73660 0 0 $X=151360 $Y=73300
X649 1336 13 12 729 1422 OR2X1 $T=157180 52780 0 180 $X=153100 $Y=46960
X650 287 13 12 64 1423 OR2X1 $T=155440 73660 0 0 $X=154840 $Y=73300
X651 1424 13 12 1425 1277 OR2X1 $T=163560 157180 1 0 $X=162960 $Y=151360
X652 313 13 12 1426 1427 OR2X1 $T=163560 157180 0 0 $X=162960 $Y=156820
X653 1340 13 12 77 1428 OR2X1 $T=184440 63220 0 180 $X=180360 $Y=57400
X654 1341 13 12 1151 324 OR2X1 $T=182120 84100 1 0 $X=181520 $Y=78280
X655 331 13 12 72 1429 OR2X1 $T=196040 63220 1 180 $X=191960 $Y=62860
X656 328 13 12 77 1430 OR2X1 $T=200100 73660 1 0 $X=199500 $Y=67840
X657 339 13 12 77 1431 OR2X1 $T=203580 42340 0 0 $X=202980 $Y=41980
X658 335 13 12 72 1432 OR2X1 $T=203580 52780 0 0 $X=202980 $Y=52420
X659 349 13 12 72 1433 OR2X1 $T=208800 31900 0 180 $X=204720 $Y=26080
X660 1162 13 12 774 1434 OR2X1 $T=214020 146740 1 0 $X=213420 $Y=140920
X661 1166 13 12 1164 1435 OR2X1 $T=215760 136300 1 0 $X=215160 $Y=130480
X662 777 13 12 769 1436 OR2X1 $T=219820 21460 1 180 $X=215740 $Y=21100
X663 1437 13 12 770 348 OR2X1 $T=222140 31900 1 180 $X=218060 $Y=31540
X664 776 13 12 768 1437 OR2X1 $T=225620 21460 1 180 $X=221540 $Y=21100
X665 365 13 12 1438 1439 OR2X1 $T=227360 125860 1 0 $X=226760 $Y=120040
X666 1440 13 12 1441 1283 OR2X1 $T=229680 146740 1 0 $X=229080 $Y=140920
X667 1346 13 12 93 1442 OR2X1 $T=238380 52780 0 180 $X=234300 $Y=46960
X668 385 13 12 79 1443 OR2X1 $T=245340 52780 0 180 $X=241260 $Y=46960
X669 1161 13 12 807 1444 OR2X1 $T=244760 146740 0 0 $X=244160 $Y=146380
X670 1445 13 12 1161 379 OR2X1 $T=250560 125860 0 180 $X=246480 $Y=120040
X671 1342 13 12 93 1446 OR2X1 $T=254040 63220 0 180 $X=249960 $Y=57400
X672 1445 13 12 1162 389 OR2X1 $T=250560 125860 1 0 $X=249960 $Y=120040
X673 1447 13 12 1448 1200 OR2X1 $T=252300 104980 1 0 $X=251700 $Y=99160
X674 797 13 12 816 1449 OR2X1 $T=256940 104980 1 180 $X=252860 $Y=104620
X675 806 13 12 811 1450 OR2X1 $T=253460 136300 0 0 $X=252860 $Y=135940
X676 1344 13 12 79 1451 OR2X1 $T=258680 63220 0 180 $X=254600 $Y=57400
X677 396 13 12 93 1452 OR2X1 $T=261580 31900 0 0 $X=260980 $Y=31540
X678 387 13 12 79 1453 OR2X1 $T=270860 31900 1 180 $X=266780 $Y=31540
X679 1189 13 12 1191 1454 OR2X1 $T=289420 21460 0 0 $X=288820 $Y=21100
X680 865 13 12 1190 1455 OR2X1 $T=295220 21460 0 0 $X=294620 $Y=21100
X681 1456 13 12 115 426 OR2X1 $T=299860 178060 1 0 $X=299260 $Y=172240
X682 1456 13 12 116 1315 OR2X1 $T=303340 178060 1 0 $X=302740 $Y=172240
X683 1348 13 12 33 1457 OR2X1 $T=310880 52780 0 180 $X=306800 $Y=46960
X684 1349 13 12 801 1458 OR2X1 $T=307980 63220 0 0 $X=307380 $Y=62860
X685 1459 13 12 1460 1292 OR2X1 $T=318420 178060 0 0 $X=317820 $Y=177700
X686 115 13 12 870 1461 OR2X1 $T=336980 178060 0 180 $X=332900 $Y=172240
X687 1210 13 12 882 1462 OR2X1 $T=341620 146740 0 0 $X=341020 $Y=146380
X688 1352 13 12 108 1463 OR2X1 $T=346840 42340 0 180 $X=342760 $Y=36520
X689 1351 13 12 108 1464 OR2X1 $T=343940 63220 0 0 $X=343340 $Y=62860
X690 1354 13 12 124 1465 OR2X1 $T=356700 63220 1 180 $X=352620 $Y=62860
X691 1353 13 12 124 1466 OR2X1 $T=357860 42340 0 0 $X=357260 $Y=41980
X692 1198 13 12 895 1467 OR2X1 $T=363660 104980 0 0 $X=363060 $Y=104620
X693 1210 13 12 886 1468 OR2X1 $T=367720 167620 0 180 $X=363640 $Y=161800
X694 899 13 12 896 479 OR2X1 $T=370620 115420 0 0 $X=370020 $Y=115060
X695 909 13 12 917 1469 OR2X1 $T=378160 146740 0 0 $X=377560 $Y=146380
X696 908 13 12 916 483 OR2X1 $T=378160 157180 1 0 $X=377560 $Y=151360
X697 1470 13 12 1210 485 OR2X1 $T=378740 115420 1 0 $X=378140 $Y=109600
X698 1470 13 12 1209 1319 OR2X1 $T=378740 125860 1 0 $X=378140 $Y=120040
X699 1209 13 12 917 1471 OR2X1 $T=381640 146740 0 0 $X=381040 $Y=146380
X700 1224 13 12 1223 1472 OR2X1 $T=382220 31900 1 0 $X=381620 $Y=26080
X701 494 13 12 137 1473 OR2X1 $T=389760 42340 1 180 $X=385680 $Y=41980
X702 1357 13 12 138 1474 OR2X1 $T=390920 63220 0 180 $X=386840 $Y=57400
X703 937 13 12 1222 1475 OR2X1 $T=388600 31900 1 0 $X=388000 $Y=26080
X704 1476 13 12 1477 1303 OR2X1 $T=392080 125860 1 180 $X=388000 $Y=125500
X705 1475 13 12 1225 493 OR2X1 $T=389760 42340 1 0 $X=389160 $Y=36520
X706 505 13 12 1478 1479 OR2X1 $T=397300 104980 1 180 $X=393220 $Y=104620
X707 514 13 12 137 1480 OR2X1 $T=409480 63220 1 180 $X=405400 $Y=62860
X708 510 13 12 137 1481 OR2X1 $T=408320 42340 0 0 $X=407720 $Y=41980
X709 1359 13 12 138 1482 OR2X1 $T=413540 63220 1 0 $X=412940 $Y=57400
X710 1358 13 12 138 1483 OR2X1 $T=415280 52780 0 0 $X=414680 $Y=52420
X711 1484 13 12 1485 978 OR2X1 $T=436160 115420 1 0 $X=435560 $Y=109600
X712 953 13 12 936 1486 OR2X1 $T=439640 21460 0 0 $X=439040 $Y=21100
X713 1487 13 12 1488 1307 OR2X1 $T=440220 167620 0 0 $X=439620 $Y=167260
X714 1489 13 12 1242 546 OR2X1 $T=444280 104980 0 180 $X=440200 $Y=99160
X715 530 13 12 151 1490 OR2X1 $T=442540 52780 0 0 $X=441940 $Y=52420
X716 952 13 12 935 1491 OR2X1 $T=448920 21460 1 180 $X=444840 $Y=21100
X717 1491 13 12 1246 548 OR2X1 $T=445440 31900 0 0 $X=444840 $Y=31540
X718 532 13 12 151 1492 OR2X1 $T=448920 73660 0 180 $X=444840 $Y=67840
X719 544 13 12 536 1251 OR2X1 $T=449500 104980 0 180 $X=445420 $Y=99160
X720 534 13 12 151 1493 OR2X1 $T=447180 84100 0 0 $X=446580 $Y=83740
X721 1494 13 12 142 1323 OR2X1 $T=451820 178060 1 180 $X=447740 $Y=177700
X722 1364 13 12 152 1495 OR2X1 $T=452400 73660 0 180 $X=448320 $Y=67840
X723 1494 13 12 144 539 OR2X1 $T=452400 178060 0 180 $X=448320 $Y=172240
X724 559 13 12 1496 1497 OR2X1 $T=454720 167620 1 180 $X=450640 $Y=167260
X725 1365 13 12 152 1498 OR2X1 $T=451820 42340 0 0 $X=451220 $Y=41980
X726 549 13 12 151 1499 OR2X1 $T=452980 31900 0 0 $X=452380 $Y=31540
X727 989 13 12 165 166 OR2X1 $T=456460 157180 1 180 $X=452380 $Y=156820
X728 1363 13 12 152 1500 OR2X1 $T=457040 73660 1 0 $X=456440 $Y=67840
X729 985 13 12 988 1501 OR2X1 $T=462260 157180 0 0 $X=461660 $Y=156820
X730 557 13 12 162 1395 OR2X1 $T=469800 104980 0 0 $X=469200 $Y=104620
X731 1374 13 12 167 1502 OR2X1 $T=472120 94540 1 0 $X=471520 $Y=88720
X732 1375 13 12 162 1503 OR2X1 $T=473280 73660 0 0 $X=472680 $Y=73300
X733 1369 13 12 167 1504 OR2X1 $T=480240 125860 0 0 $X=479640 $Y=125500
X734 1371 13 12 167 1505 OR2X1 $T=484880 31900 1 0 $X=484280 $Y=26080
X735 1377 13 12 162 1506 OR2X1 $T=488940 31900 0 0 $X=488340 $Y=31540
X736 1507 13 12 1508 1040 OR2X1 $T=492420 104980 0 180 $X=488340 $Y=99160
X737 1378 13 12 162 1509 OR2X1 $T=489520 52780 1 0 $X=488920 $Y=46960
X738 1372 13 12 167 1510 OR2X1 $T=489520 63220 1 0 $X=488920 $Y=57400
X739 1376 13 12 162 1511 OR2X1 $T=489520 94540 0 0 $X=488920 $Y=94180
X740 1373 13 12 167 1512 OR2X1 $T=490100 73660 0 0 $X=489500 $Y=73300
X741 1379 13 12 183 573 OR2X1 $T=498220 136300 1 0 $X=497620 $Y=130480
X742 563 13 12 183 1513 OR2X1 $T=501120 42340 0 0 $X=500520 $Y=41980
X743 570 13 12 183 1514 OR2X1 $T=505760 84100 1 0 $X=505160 $Y=78280
X744 1260 13 12 1262 563 OR2X1 $T=510400 31900 0 180 $X=506320 $Y=26080
X745 1513 13 12 1058 1515 OR2X1 $T=507500 52780 0 0 $X=506900 $Y=52420
X746 566 13 12 183 1516 OR2X1 $T=509820 94540 0 0 $X=509220 $Y=94180
X747 1381 13 12 1035 585 OR2X1 $T=511560 115420 0 0 $X=510960 $Y=115060
X748 585 13 12 186 577 OR2X1 $T=515040 125860 1 180 $X=510960 $Y=125500
X749 1380 13 12 186 1517 OR2X1 $T=513300 94540 0 0 $X=512700 $Y=94180
X750 1075 13 12 1261 1518 OR2X1 $T=517360 31900 1 180 $X=513280 $Y=31540
X751 1518 13 12 186 1519 OR2X1 $T=516780 42340 1 0 $X=516180 $Y=36520
X752 1382 13 12 186 1520 OR2X1 $T=520260 84100 1 180 $X=516180 $Y=83740
X753 1519 13 12 1057 1521 OR2X1 $T=519100 52780 0 0 $X=518500 $Y=52420
X754 1324 649 13 12 638 NOR2BXL $T=50460 94540 0 0 $X=49860 $Y=94180
X755 1325 650 13 12 637 NOR2BXL $T=51620 94540 1 0 $X=51020 $Y=88720
X756 1522 657 13 12 1523 NOR2BXL $T=62640 73660 0 180 $X=58560 $Y=67840
X757 1524 1525 13 12 657 NOR2BXL $T=67280 73660 0 180 $X=63200 $Y=67840
X758 236 647 13 12 663 NOR2BXL $T=67860 42340 0 180 $X=63780 $Y=36520
X759 232 1097 13 12 234 NOR2BXL $T=67860 125860 0 180 $X=63780 $Y=120040
X760 1399 31 13 12 230 NOR2BXL $T=70180 52780 0 0 $X=69580 $Y=52420
X761 1400 1389 13 12 1094 NOR2BXL $T=77720 115420 1 180 $X=73640 $Y=115060
X762 251 677 13 12 599 NOR2BXL $T=88160 52780 0 180 $X=84080 $Y=46960
X763 248 43 13 12 41 NOR2BXL $T=96280 188500 1 0 $X=95680 $Y=182680
X764 269 42 13 12 29 NOR2BXL $T=106140 178060 1 180 $X=102060 $Y=177700
X765 260 1332 13 12 48 NOR2BXL $T=114840 104980 1 0 $X=114240 $Y=99160
X766 278 710 13 12 1127 NOR2BXL $T=132820 157180 1 180 $X=128740 $Y=156820
X767 1412 41 13 12 62 NOR2BXL $T=138040 188500 0 180 $X=133960 $Y=182680
X768 1526 49 13 12 1414 NOR2BXL $T=151960 157180 0 0 $X=151360 $Y=156820
X769 285 307 13 12 1136 NOR2BXL $T=156600 104980 0 180 $X=152520 $Y=99160
X770 309 303 13 12 801 NOR2BXL $T=153120 167620 1 0 $X=152520 $Y=161800
X771 1527 324 13 12 72 NOR2BXL $T=186180 84100 1 180 $X=182100 $Y=83740
X772 1528 72 13 12 337 NOR2BXL $T=196040 84100 1 180 $X=191960 $Y=83740
X773 1529 1161 13 12 1435 NOR2BXL $T=214020 146740 0 180 $X=209940 $Y=140920
X774 339 1436 13 12 770 NOR2BXL $T=215180 31900 0 0 $X=214580 $Y=31540
X775 359 796 13 12 1166 NOR2BXL $T=231420 115420 1 0 $X=230820 $Y=109600
X776 377 371 13 12 33 NOR2BXL $T=236060 115420 1 180 $X=231980 $Y=115060
X777 1530 1345 13 12 779 NOR2BXL $T=241280 73660 1 180 $X=237200 $Y=73300
X778 1445 807 13 12 811 NOR2BXL $T=249980 136300 0 0 $X=249380 $Y=135940
X779 1531 613 13 12 807 NOR2BXL $T=268540 136300 0 180 $X=264460 $Y=130480
X780 1532 806 13 12 613 NOR2BXL $T=272020 136300 1 0 $X=271420 $Y=130480
X781 1533 33 13 12 416 NOR2BXL $T=281300 73660 0 0 $X=280700 $Y=73300
X782 1456 96 13 12 1179 NOR2BXL $T=294640 178060 0 180 $X=290560 $Y=172240
X783 1534 1350 13 12 826 NOR2BXL $T=302760 73660 0 180 $X=298680 $Y=67840
X784 1312 115 13 12 848 NOR2BXL $T=310300 178060 0 180 $X=306220 $Y=172240
X785 456 116 13 12 871 NOR2BXL $T=341620 178060 0 180 $X=337540 $Y=172240
X786 1535 891 13 12 863 NOR2BXL $T=345100 31900 0 180 $X=341020 $Y=26080
X787 1536 1355 13 12 1208 NOR2BXL $T=350900 84100 0 180 $X=346820 $Y=78280
X788 1537 1209 13 12 883 NOR2BXL $T=356120 167620 0 180 $X=352040 $Y=161800
X789 1538 906 13 12 909 NOR2BXL $T=370620 146740 0 180 $X=366540 $Y=140920
X790 1539 621 13 12 864 NOR2BXL $T=368880 21460 0 0 $X=368280 $Y=21100
X791 1540 908 13 12 906 NOR2BXL $T=374100 146740 0 180 $X=370020 $Y=140920
X792 1318 1210 13 12 860 NOR2BXL $T=381640 115420 1 180 $X=377560 $Y=115060
X793 487 1209 13 12 1469 NOR2BXL $T=381640 136300 0 180 $X=377560 $Y=130480
X794 1470 1199 13 12 1201 NOR2BXL $T=379320 104980 0 0 $X=378720 $Y=104620
X795 1357 1472 13 12 1225 NOR2BXL $T=383960 42340 1 0 $X=383360 $Y=36520
X796 1541 490 13 12 1542 NOR2BXL $T=406580 125860 0 180 $X=402500 $Y=120040
X797 1543 137 13 12 507 NOR2BXL $T=410060 84100 0 180 $X=405980 $Y=78280
X798 1544 1360 13 12 923 NOR2BXL $T=419340 84100 1 0 $X=418740 $Y=78280
X799 1322 144 13 12 945 NOR2BXL $T=437900 178060 0 180 $X=433820 $Y=172240
X800 1365 1486 13 12 1246 NOR2BXL $T=440800 31900 0 0 $X=440200 $Y=31540
X801 1494 986 13 12 948 NOR2BXL $T=452400 178060 1 0 $X=451800 $Y=172240
X802 553 1366 13 12 151 NOR2BXL $T=455880 84100 0 0 $X=455280 $Y=83740
X803 1545 622 13 12 165 NOR2BXL $T=461680 157180 1 180 $X=457600 $Y=156820
X804 1546 168 13 12 622 NOR2BXL $T=472120 157180 1 180 $X=468040 $Y=156820
X805 1547 991 13 12 981 NOR2BXL $T=473860 21460 1 180 $X=469780 $Y=21100
X806 1548 992 13 12 980 NOR2BXL $T=479660 21460 1 180 $X=475580 $Y=21100
X807 639 224 13 12 643 1549 OA21X1 $T=50460 136300 1 0 $X=49860 $Y=130480
X808 651 1549 13 12 23 1550 OA21X1 $T=53360 136300 0 0 $X=52760 $Y=135940
X809 654 237 13 12 658 1525 OA21X1 $T=57420 52780 0 0 $X=56820 $Y=52420
X810 664 1522 13 12 667 1327 OA21X1 $T=63800 94540 0 180 $X=57980 $Y=88720
X811 674 1401 13 12 31 1551 OA21X1 $T=70180 136300 0 0 $X=69580 $Y=135940
X812 665 1524 13 12 668 1398 OA21X1 $T=73080 94540 0 0 $X=72480 $Y=94180
X813 1112 1329 13 12 1115 258 OA21X1 $T=114840 63220 1 180 $X=109020 $Y=62860
X814 1113 1331 13 12 1116 262 OA21X1 $T=120640 63220 1 180 $X=114820 $Y=62860
X815 1552 1384 13 12 309 1420 OA21X1 $T=133980 167620 1 0 $X=133380 $Y=161800
X816 53 269 13 12 284 289 OA21X1 $T=138620 178060 0 0 $X=138020 $Y=177700
X817 711 53 13 12 1553 1554 OA21X1 $T=139200 167620 1 0 $X=138600 $Y=161800
X818 30 53 13 12 289 1553 OA21X1 $T=139780 178060 1 0 $X=139180 $Y=172240
X819 53 278 13 12 1553 1555 OA21X1 $T=140360 157180 0 0 $X=139760 $Y=156820
X820 1132 53 13 12 1555 1556 OA21X1 $T=140940 157180 1 0 $X=140340 $Y=151360
X821 291 1554 13 12 33 1419 OA21X1 $T=144420 167620 1 0 $X=143820 $Y=161800
X822 740 1337 13 12 1139 293 OA21X1 $T=150220 52780 1 180 $X=144400 $Y=52420
X823 1144 1557 13 12 64 1558 OA21X1 $T=150220 115420 1 0 $X=149620 $Y=109600
X824 736 734 13 12 1147 1335 OA21X1 $T=160080 31900 1 180 $X=154260 $Y=31540
X825 735 733 13 12 1146 1336 OA21X1 $T=164140 42340 0 180 $X=158320 $Y=36520
X826 1164 1162 13 12 1559 1560 OA21X1 $T=219820 125860 0 0 $X=219220 $Y=125500
X827 1162 359 13 12 1561 1559 OA21X1 $T=227360 115420 0 0 $X=226760 $Y=115060
X828 1562 1386 13 12 377 1448 OA21X1 $T=234900 115420 1 0 $X=234300 $Y=109600
X829 373 1563 13 12 801 1447 OA21X1 $T=247080 104980 1 0 $X=246480 $Y=99160
X830 797 1162 13 12 1561 1563 OA21X1 $T=252300 104980 1 180 $X=246480 $Y=104620
X831 615 1181 13 12 808 395 OA21X1 $T=254040 31900 1 0 $X=253440 $Y=26080
X832 857 1455 13 12 830 428 OA21X1 $T=309140 31900 0 180 $X=303320 $Y=26080
X833 858 1454 13 12 831 434 OA21X1 $T=313780 31900 1 180 $X=307960 $Y=31540
X834 883 1210 13 12 1564 1565 OA21X1 $T=347420 167620 1 0 $X=346820 $Y=161800
X835 1209 480 13 12 488 489 OA21X1 $T=381640 125860 0 0 $X=381040 $Y=125500
X836 1209 484 13 12 1566 1567 OA21X1 $T=385120 146740 0 0 $X=384520 $Y=146380
X837 899 1209 13 12 1567 499 OA21X1 $T=392660 136300 1 0 $X=392060 $Y=130480
X838 1239 546 13 12 151 1484 OA21X1 $T=439640 104980 0 180 $X=433820 $Y=99160
X839 550 142 13 12 164 541 OA21X1 $T=451820 188500 0 180 $X=446000 $Y=182680
X840 1255 1370 13 12 162 1507 OA21X1 $T=490100 104980 0 0 $X=489500 $Y=104620
X841 1032 577 13 12 573 579 OA21X1 $T=506340 136300 1 0 $X=505740 $Y=130480
X842 1263 1568 13 12 189 1569 OA21X1 $T=517940 146740 0 0 $X=517340 $Y=146380
X843 1326 227 13 12 23 223 MXI2XL $T=56260 115420 0 180 $X=51020 $Y=109600
X844 32 1273 13 12 33 242 MXI2XL $T=71340 167620 1 180 $X=66100 $Y=167260
X845 1522 240 13 12 31 1524 MXI2XL $T=70760 73660 1 0 $X=70160 $Y=67840
X846 252 1114 13 12 40 244 MXI2XL $T=88740 63220 0 180 $X=83500 $Y=57400
X847 1570 1274 13 12 33 1571 MXI2XL $T=101500 167620 1 0 $X=100900 $Y=161800
X848 1331 271 13 12 48 1329 MXI2XL $T=114260 63220 0 180 $X=109020 $Y=57400
X849 1572 1276 13 12 33 297 MXI2XL $T=148480 136300 0 180 $X=143240 $Y=130480
X850 57 65 13 12 33 61 MXI2XL $T=144420 188500 1 0 $X=143820 $Y=182680
X851 1337 316 13 12 729 299 MXI2XL $T=154280 52780 0 0 $X=153680 $Y=52420
X852 323 1278 13 12 33 1573 MXI2XL $T=183860 136300 1 0 $X=183260 $Y=130480
X853 78 1279 13 12 33 1574 MXI2XL $T=189660 178060 0 180 $X=184420 $Y=172240
X854 1575 346 13 12 72 1576 MXI2XL $T=204740 52780 0 180 $X=199500 $Y=46960
X855 341 1282 13 12 33 334 MXI2XL $T=209380 157180 0 180 $X=204140 $Y=151360
X856 351 1281 13 12 33 357 MXI2XL $T=214020 115420 1 0 $X=213420 $Y=109600
X857 353 1280 13 12 33 1577 MXI2XL $T=219820 125860 1 180 $X=214580 $Y=125500
X858 1578 1284 13 12 33 384 MXI2XL $T=244180 136300 1 180 $X=238940 $Y=135940
X859 397 407 13 12 93 392 MXI2XL $T=261000 42340 1 180 $X=255760 $Y=41980
X860 413 1285 13 12 108 410 MXI2XL $T=280140 167620 0 180 $X=274900 $Y=161800
X861 403 1286 13 12 33 415 MXI2XL $T=277820 94540 0 0 $X=277220 $Y=94180
X862 1579 1290 13 12 108 110 MXI2XL $T=277820 188500 1 0 $X=277220 $Y=182680
X863 422 1289 13 12 33 1580 MXI2XL $T=298700 115420 1 180 $X=293460 $Y=115060
X864 428 444 13 12 801 434 MXI2XL $T=306820 42340 1 0 $X=306220 $Y=36520
X865 1581 1293 13 12 108 1582 MXI2XL $T=315520 157180 1 180 $X=310280 $Y=156820
X866 1454 1213 13 12 33 1455 MXI2XL $T=317840 31900 0 180 $X=312600 $Y=26080
X867 448 1294 13 12 108 451 MXI2XL $T=335820 104980 0 180 $X=330580 $Y=99160
X868 1583 1299 13 12 108 1584 MXI2XL $T=335240 125860 0 0 $X=334640 $Y=125500
X869 1585 1295 13 12 108 1586 MXI2XL $T=335240 157180 1 0 $X=334640 $Y=151360
X870 1564 1296 13 12 108 1587 MXI2XL $T=348000 157180 1 180 $X=342760 $Y=156820
X871 1535 462 13 12 108 1539 MXI2XL $T=350320 31900 1 180 $X=345080 $Y=31540
X872 1588 464 13 12 108 1589 MXI2XL $T=350320 31900 0 0 $X=349720 $Y=31540
X873 455 1298 13 12 108 1590 MXI2XL $T=350320 84100 0 0 $X=349720 $Y=83740
X874 1591 1301 13 12 108 470 MXI2XL $T=370620 104980 0 0 $X=370020 $Y=104620
X875 1592 1302 13 12 108 1566 MXI2XL $T=390340 157180 1 180 $X=385100 $Y=156820
X876 523 1306 13 12 137 528 MXI2XL $T=422820 157180 0 0 $X=422220 $Y=156820
X877 537 1308 13 12 137 1593 MXI2XL $T=444860 146740 0 180 $X=439620 $Y=140920
X878 1594 1310 13 12 137 1595 MXI2XL $T=473860 125860 0 0 $X=473260 $Y=125500
X879 1548 567 13 12 167 1547 MXI2XL $T=486040 21460 0 0 $X=485440 $Y=21100
X880 581 191 13 12 151 188 MXI2XL $T=512720 188500 0 180 $X=507480 $Y=182680
X881 197 196 13 12 151 588 MXI2XL $T=524900 188500 0 180 $X=519660 $Y=182680
X882 254 1110 13 12 698 1403 AND3X1 $T=85260 94540 1 180 $X=80020 $Y=94180
X883 246 686 13 12 1103 1596 AND3X1 $T=91640 115420 0 0 $X=91040 $Y=115060
X884 258 1117 13 12 712 1405 AND3X1 $T=110200 84100 0 0 $X=109600 $Y=83740
X885 262 1118 13 12 713 1333 AND3X1 $T=116580 84100 0 0 $X=115980 $Y=83740
X886 293 1133 13 12 717 1417 AND3X1 $T=144420 73660 0 180 $X=139180 $Y=67840
X887 288 1134 13 12 718 1338 AND3X1 $T=146740 73660 0 0 $X=146140 $Y=73300
X888 329 1148 13 12 737 1340 AND3X1 $T=189080 63220 0 180 $X=183840 $Y=57400
X889 332 745 13 12 748 326 AND3X1 $T=187340 73660 0 0 $X=186740 $Y=73300
X890 326 751 13 12 1151 337 AND3X1 $T=187920 84100 0 0 $X=187320 $Y=83740
X891 325 632 13 12 1158 1597 AND3X1 $T=190240 94540 1 0 $X=189640 $Y=88720
X892 340 1155 13 12 757 1576 AND3X1 $T=196040 42340 1 180 $X=190800 $Y=41980
X893 336 1149 13 12 738 331 AND3X1 $T=196040 63220 0 180 $X=190800 $Y=57400
X894 348 1154 13 12 756 1575 AND3X1 $T=204160 42340 0 180 $X=198920 $Y=36520
X895 388 788 13 12 791 385 AND3X1 $T=245920 42340 0 180 $X=240680 $Y=36520
X896 1530 631 13 12 1168 1598 AND3X1 $T=248240 84100 0 180 $X=243000 $Y=78280
X897 386 1173 13 12 1175 391 AND3X1 $T=249400 52780 1 0 $X=248800 $Y=46960
X898 395 787 13 12 790 1346 AND3X1 $T=254620 42340 0 180 $X=249380 $Y=36520
X899 1536 616 13 12 1221 1599 AND3X1 $T=356700 84100 0 0 $X=356100 $Y=83740
X900 493 1227 13 12 1229 509 AND3X1 $T=397880 52780 1 0 $X=397280 $Y=46960
X901 513 919 13 12 913 517 AND3X1 $T=403100 73660 0 180 $X=397860 $Y=67840
X902 517 1232 13 12 922 507 AND3X1 $T=401360 84100 1 0 $X=400760 $Y=78280
X903 509 925 13 12 932 513 AND3X1 $T=405420 52780 0 0 $X=404820 $Y=52420
X904 1544 1233 13 12 1235 1600 AND3X1 $T=415860 84100 1 180 $X=410620 $Y=83740
X905 531 963 13 12 969 533 AND3X1 $T=440800 73660 0 180 $X=435560 $Y=67840
X906 533 972 13 12 975 1601 AND3X1 $T=441380 94540 0 180 $X=436140 $Y=88720
X907 548 960 13 12 966 529 AND3X1 $T=444280 42340 1 180 $X=439040 $Y=41980
X908 529 957 13 12 954 531 AND3X1 $T=440220 63220 1 0 $X=439620 $Y=57400
X909 553 976 13 12 973 544 AND3X1 $T=455300 84100 1 180 $X=450060 $Y=83740
X910 569 1053 13 12 1050 565 AND3X1 $T=504600 84100 0 180 $X=499360 $Y=78280
X911 565 1060 13 12 1047 575 AND3X1 $T=502860 104980 0 0 $X=502260 $Y=104620
X912 586 1033 13 12 1030 1602 AND3X1 $T=516780 136300 1 180 $X=511540 $Y=135940
X913 57 13 12 1409 49 54 41 33 AOI221XL $T=127600 188500 0 180 $X=121200 $Y=182680
X914 53 13 12 732 1556 1603 1416 1526 AOI221XL $T=147900 146740 0 0 $X=147300 $Y=146380
X915 1560 13 12 1434 1162 1604 774 1529 AOI221XL $T=223300 146740 0 180 $X=216900 $Y=140920
X916 1161 13 12 807 384 1605 1444 801 AOI221XL $T=249980 136300 1 180 $X=243580 $Y=135940
X917 93 13 12 800 79 405 1181 1606 AOI221XL $T=253460 31900 0 180 $X=247060 $Y=26080
X918 801 13 12 833 33 436 834 444 AOI221XL $T=313780 42340 1 0 $X=313180 $Y=36520
X919 1210 13 12 886 1565 1592 1468 1537 AOI221XL $T=361920 167620 0 180 $X=355520 $Y=161800
X920 124 13 12 1216 108 468 1217 465 AOI221XL $T=367140 42340 1 0 $X=366540 $Y=36520
X921 1566 13 12 1471 1209 1607 917 124 AOI221XL $T=384540 157180 1 180 $X=378140 $Y=156820
X922 1397 645 13 12 646 1396 642 662 BMXIX2 $T=49880 104980 1 180 $X=34200 $Y=104620
X923 1325 641 13 12 642 1324 653 669 BMXIX2 $T=50460 94540 1 180 $X=34780 $Y=94180
X924 649 653 13 12 23 650 638 666 BMXIX2 $T=39440 84100 0 0 $X=38840 $Y=83740
X925 226 651 13 12 652 1549 653 676 BMXIX2 $T=55100 146740 0 180 $X=39420 $Y=140920
X926 229 654 13 12 655 237 672 600 BMXIX2 $T=53360 42340 0 0 $X=52760 $Y=41980
X927 233 674 13 12 675 1401 672 682 BMXIX2 $T=67280 136300 1 0 $X=66680 $Y=130480
X928 1327 660 13 12 661 1398 672 699 BMXIX2 $T=69020 104980 1 0 $X=68420 $Y=99160
X929 235 1096 13 12 1097 1400 672 687 BMXIX2 $T=69600 125860 1 0 $X=69000 $Y=120040
X930 247 1102 13 12 1103 1403 40 702 BMXIX2 $T=74240 104980 0 0 $X=73640 $Y=104620
X931 1402 1109 13 12 1110 253 40 714 BMXIX2 $T=84100 84100 0 0 $X=83500 $Y=83740
X932 263 1117 13 12 1118 259 705 719 BMXIX2 $T=109620 73660 0 0 $X=109020 $Y=73300
X933 1405 1120 13 12 1121 1333 48 728 BMXIX2 $T=109620 94540 1 0 $X=109020 $Y=88720
X934 1330 692 13 12 693 1328 705 725 BMXIX2 $T=110780 42340 0 0 $X=110180 $Y=41980
X935 1406 694 13 12 695 1407 692 742 BMXIX2 $T=110780 52780 0 0 $X=110180 $Y=52420
X936 1410 712 13 12 713 1408 1118 722 BMXIX2 $T=126440 84100 0 180 $X=110760 $Y=78280
X937 1335 1128 13 12 1129 1336 729 758 BMXIX2 $T=141520 42340 1 0 $X=140920 $Y=36520
X938 287 1133 13 12 1134 294 729 739 BMXIX2 $T=141520 63220 0 0 $X=140920 $Y=62860
X939 1338 720 13 12 721 1417 729 750 BMXIX2 $T=145000 84100 1 0 $X=144400 $Y=78280
X940 286 1144 13 12 1145 1557 729 755 BMXIX2 $T=146160 104980 0 0 $X=145560 $Y=104620
X941 1413 723 13 12 724 1422 1128 761 BMXIX2 $T=146740 42340 0 0 $X=146140 $Y=41980
X942 1423 717 13 12 718 1421 1134 747 BMXIX2 $T=147320 73660 1 0 $X=146720 $Y=67840
X943 1383 305 13 12 306 1608 801 71 BMXIX2 $T=151380 178060 1 0 $X=150780 $Y=172240
X944 1339 1141 13 12 1142 301 726 752 BMXIX2 $T=155440 94540 1 0 $X=154840 $Y=88720
X945 1341 1151 13 12 1152 327 72 780 BMXIX2 $T=180960 84100 0 180 $X=165280 $Y=78280
X946 1428 748 13 12 749 1429 746 783 BMXIX2 $T=177480 63220 0 0 $X=176880 $Y=62860
X947 1340 745 13 12 746 331 72 786 BMXIX2 $T=180960 73660 1 0 $X=180360 $Y=67840
X948 1431 756 13 12 757 1433 1155 792 BMXIX2 $T=198360 31900 0 0 $X=197760 $Y=31540
X949 328 1148 13 12 1149 335 72 821 BMXIX2 $T=198940 63220 0 0 $X=198340 $Y=62860
X950 1430 737 13 12 738 1432 1148 824 BMXIX2 $T=200100 63220 1 0 $X=199500 $Y=57400
X951 90 91 13 12 89 92 79 798 BMXIX2 $T=210540 188500 1 0 $X=209940 $Y=182680
X952 1436 770 13 12 771 1437 72 810 BMXIX2 $T=211120 31900 1 0 $X=210520 $Y=26080
X953 339 1154 13 12 1155 349 72 789 BMXIX2 $T=211700 42340 0 0 $X=211100 $Y=41980
X954 1346 1173 13 12 1174 385 79 835 BMXIX2 $T=233740 42340 0 0 $X=233140 $Y=41980
X955 1342 784 13 12 785 1344 79 841 BMXIX2 $T=233740 63220 1 0 $X=233140 $Y=57400
X956 369 778 13 12 779 1345 79 853 BMXIX2 $T=234320 73660 1 0 $X=233720 $Y=67840
X957 1442 1175 13 12 1176 1443 1174 838 BMXIX2 $T=234900 52780 0 0 $X=234300 $Y=52420
X958 1385 381 13 12 382 1609 33 897 BMXIX2 $T=241860 115420 1 0 $X=241260 $Y=109600
X959 1452 790 13 12 791 1453 787 832 BMXIX2 $T=242440 31900 0 0 $X=241840 $Y=31540
X960 1446 781 13 12 782 1451 784 827 BMXIX2 $T=245340 63220 0 0 $X=244740 $Y=62860
X961 396 787 13 12 788 387 79 859 BMXIX2 $T=256360 42340 1 0 $X=255760 $Y=36520
X962 418 825 13 12 826 1350 801 875 BMXIX2 $T=288840 63220 0 0 $X=288240 $Y=62860
X963 1347 1187 13 12 1188 432 851 617 BMXIX2 $T=295800 73660 0 0 $X=295200 $Y=73300
X964 1348 1194 13 12 1195 1349 801 878 BMXIX2 $T=301600 52780 0 0 $X=301000 $Y=52420
X965 1457 839 13 12 840 1458 1194 881 BMXIX2 $T=302180 63220 1 0 $X=301580 $Y=57400
X966 1352 1204 13 12 1205 1353 124 927 BMXIX2 $T=339880 52780 1 0 $X=339280 $Y=46960
X967 458 1207 13 12 1208 1355 124 924 BMXIX2 $T=341620 73660 0 0 $X=341020 $Y=73300
X968 1351 879 13 12 880 1354 124 921 BMXIX2 $T=342200 63220 1 0 $X=341600 $Y=57400
X969 1463 876 13 12 877 1466 1204 934 BMXIX2 $T=342780 42340 0 0 $X=342180 $Y=41980
X970 1464 873 13 12 874 1465 879 915 BMXIX2 $T=343360 73660 1 0 $X=342760 $Y=67840
X971 1474 1229 13 12 1230 1473 1228 959 BMXIX2 $T=381640 52780 0 0 $X=381040 $Y=52420
X972 1357 1227 13 12 1228 494 137 968 BMXIX2 $T=382800 52780 1 0 $X=382200 $Y=46960
X973 1472 1225 13 12 1226 1475 137 962 BMXIX2 $T=383960 31900 0 0 $X=383360 $Y=31540
X974 1387 511 13 12 512 1610 108 990 BMXIX2 $T=397880 136300 0 0 $X=397280 $Y=135940
X975 1611 521 13 12 522 1362 124 950 BMXIX2 $T=402520 115420 1 0 $X=401920 $Y=109600
X976 1541 515 13 12 516 1612 124 987 BMXIX2 $T=406580 125860 1 0 $X=405980 $Y=120040
X977 510 925 13 12 926 1358 138 956 BMXIX2 $T=407740 52780 1 0 $X=407140 $Y=46960
X978 1480 913 13 12 914 1482 919 977 BMXIX2 $T=407740 73660 1 0 $X=407140 $Y=67840
X979 518 922 13 12 923 1360 138 974 BMXIX2 $T=408900 73660 0 0 $X=408300 $Y=73300
X980 514 919 13 12 920 1359 138 971 BMXIX2 $T=409480 63220 0 0 $X=408880 $Y=62860
X981 1481 932 13 12 933 1483 925 965 BMXIX2 $T=411800 42340 0 0 $X=411200 $Y=41980
X982 1486 1246 13 12 1247 1491 151 995 BMXIX2 $T=438480 31900 1 0 $X=437880 $Y=26080
X983 1365 960 13 12 961 549 151 998 BMXIX2 $T=444280 42340 1 0 $X=443680 $Y=36520
X984 535 1244 13 12 1245 545 1242 1022 BMXIX2 $T=444280 94540 0 0 $X=443680 $Y=94180
X985 1498 966 13 12 967 1499 961 1001 BMXIX2 $T=444860 52780 1 0 $X=444260 $Y=46960
X986 534 975 13 12 976 1366 152 1025 BMXIX2 $T=445440 84100 1 0 $X=444840 $Y=78280
X987 1363 957 13 12 958 530 151 1004 BMXIX2 $T=446020 52780 0 0 $X=445420 $Y=52420
X988 1492 969 13 12 970 1495 963 1013 BMXIX2 $T=446020 73660 0 0 $X=445420 $Y=73300
X989 1490 954 13 12 955 1500 957 1007 BMXIX2 $T=447180 63220 1 0 $X=446580 $Y=57400
X990 532 963 13 12 964 1364 152 1010 BMXIX2 $T=448340 63220 0 0 $X=447740 $Y=62860
X991 1493 972 13 12 973 554 975 1016 BMXIX2 $T=450660 94540 1 0 $X=450060 $Y=88720
X992 1511 1014 13 12 1015 1502 1023 1037 BMXIX2 $T=483140 84100 1 180 $X=467460 $Y=83740
X993 1368 561 13 12 562 1613 137 1028 BMXIX2 $T=470960 178060 1 0 $X=470360 $Y=172240
X994 1395 1020 13 12 1021 1504 1249 1031 BMXIX2 $T=472700 115420 0 0 $X=472100 $Y=115060
X995 557 1249 13 12 1250 1369 167 1034 BMXIX2 $T=473860 125860 1 0 $X=473260 $Y=120040
X996 1505 999 13 12 1000 1506 997 1043 BMXIX2 $T=478500 42340 0 0 $X=477900 $Y=41980
X997 1509 1005 13 12 1006 1510 1002 1055 BMXIX2 $T=494160 63220 1 180 $X=478480 $Y=62860
X998 1376 1023 13 12 1024 1374 167 1049 BMXIX2 $T=480820 94540 1 0 $X=480220 $Y=88720
X999 1371 996 13 12 997 1377 162 1059 BMXIX2 $T=484880 42340 1 0 $X=484280 $Y=36520
X1000 1378 1002 13 12 1003 1372 167 1046 BMXIX2 $T=484880 52780 0 0 $X=484280 $Y=52420
X1001 1375 1008 13 12 1009 1373 167 1052 BMXIX2 $T=484880 73660 1 0 $X=484280 $Y=67840
X1002 1503 1011 13 12 1012 1512 1008 1062 BMXIX2 $T=484880 84100 1 0 $X=484280 $Y=78280
X1003 566 1060 13 12 1061 1380 186 1087 BMXIX2 $T=504020 94540 1 0 $X=503420 $Y=88720
X1004 563 1057 13 12 1058 1518 186 1090 BMXIX2 $T=504600 42340 0 0 $X=504000 $Y=41980
X1005 570 1053 13 12 1054 1382 186 1081 BMXIX2 $T=505760 73660 1 0 $X=505160 $Y=67840
X1006 576 1035 13 12 1036 1381 186 1067 BMXIX2 $T=506920 115420 1 0 $X=506320 $Y=109600
X1007 1513 1041 13 12 1042 1519 1057 1093 BMXIX2 $T=509820 52780 1 0 $X=509220 $Y=46960
X1008 1515 1044 13 12 1045 1521 1041 1078 BMXIX2 $T=509820 63220 1 0 $X=509220 $Y=57400
X1009 1514 1050 13 12 1051 1520 1053 1084 BMXIX2 $T=510400 84100 1 0 $X=509800 $Y=78280
X1010 1516 1047 13 12 1048 1517 1060 1070 BMXIX2 $T=510980 104980 1 0 $X=510380 $Y=99160
X1011 267 691 13 12 703 276 ADDHX1 $T=128760 42340 1 0 $X=128160 $Y=36520
X1012 1552 710 13 12 53 305 ADDHX1 $T=131660 167620 0 0 $X=131060 $Y=167260
X1013 1391 1127 13 12 49 367 ADDHX1 $T=160080 167620 0 0 $X=159480 $Y=167260
X1014 1426 1131 13 12 53 355 ADDHX1 $T=167040 167620 1 0 $X=166440 $Y=161800
X1015 1438 1163 13 12 1162 430 ADDHX1 $T=225040 125860 0 0 $X=224440 $Y=125500
X1016 1562 796 13 12 1162 381 ADDHX1 $T=232580 104980 0 0 $X=231980 $Y=104620
X1017 1393 1166 13 12 1161 424 ADDHX1 $T=237800 125860 1 0 $X=237200 $Y=120040
X1018 1606 1182 13 12 615 393 ADDHX1 $T=247660 21460 1 0 $X=247060 $Y=15640
X1019 119 1179 13 12 115 113 ADDHX1 $T=302760 188500 0 180 $X=292880 $Y=182680
X1020 1478 1201 13 12 1210 521 ADDHX1 $T=389760 115420 1 0 $X=389160 $Y=109600
X1021 503 895 13 12 1210 511 ADDHX1 $T=397880 136300 1 0 $X=397280 $Y=130480
X1022 1361 1199 13 12 1209 515 ADDHX1 $T=407740 115420 0 0 $X=407140 $Y=115060
X1023 1496 948 13 12 144 561 ADDHX1 $T=455880 167620 0 0 $X=455280 $Y=167260
X1024 1614 988 13 12 144 176 ADDHX1 $T=469800 188500 1 0 $X=469200 $Y=182680
X1025 1367 986 13 12 142 178 ADDHX1 $T=472700 178060 0 0 $X=472100 $Y=177700
X1026 639 13 12 1326 643 225 AO21X1 $T=56840 136300 1 0 $X=56240 $Y=130480
X1027 654 13 12 230 658 1523 AO21X1 $T=64960 63220 0 180 $X=59140 $Y=57400
X1028 651 13 12 225 1550 673 AO21X1 $T=61480 136300 0 0 $X=60880 $Y=135940
X1029 674 13 12 232 1551 681 AO21X1 $T=75400 136300 0 0 $X=74800 $Y=135940
X1030 628 13 12 1596 680 1615 AO21X1 $T=96280 115420 0 0 $X=95680 $Y=115060
X1031 703 13 12 690 688 1328 AO21X1 $T=104400 31900 1 180 $X=98580 $Y=31540
X1032 691 13 12 704 689 1330 AO21X1 $T=116580 42340 0 180 $X=110760 $Y=36520
X1033 627 13 12 265 705 1616 AO21X1 $T=124120 115420 1 0 $X=123520 $Y=109600
X1034 33 13 12 58 54 60 AO21X1 $T=127600 188500 1 0 $X=127000 $Y=182680
X1035 53 13 12 707 280 1384 AO21X1 $T=128180 178060 1 0 $X=127580 $Y=172240
X1036 53 13 12 270 275 280 AO21X1 $T=128180 178060 0 0 $X=127580 $Y=177700
X1037 53 13 12 279 1384 313 AO21X1 $T=135140 157180 0 0 $X=134540 $Y=156820
X1038 53 13 12 1415 296 291 AO21X1 $T=150800 167620 1 180 $X=144980 $Y=167260
X1039 49 13 12 1415 283 303 AO21X1 $T=150800 167620 0 0 $X=150200 $Y=167260
X1040 740 13 12 300 1139 287 AO21X1 $T=151380 63220 1 0 $X=150780 $Y=57400
X1041 295 13 12 290 801 1617 AO21X1 $T=151380 178060 0 0 $X=150780 $Y=177700
X1042 292 13 12 1603 801 1618 AO21X1 $T=153700 146740 0 0 $X=153100 $Y=146380
X1043 1144 13 12 285 1558 744 AO21X1 $T=157180 115420 1 0 $X=156580 $Y=109600
X1044 754 13 12 1597 77 1619 AO21X1 $T=190240 94540 0 0 $X=189640 $Y=94180
X1045 760 13 12 1576 1160 328 AO21X1 $T=196040 52780 1 180 $X=190220 $Y=52420
X1046 759 13 12 1575 1159 335 AO21X1 $T=198360 52780 0 0 $X=197760 $Y=52420
X1047 632 13 12 1527 1528 1169 AO21X1 $T=199520 84100 0 0 $X=198920 $Y=83740
X1048 1162 13 12 360 1386 365 AO21X1 $T=222140 115420 0 0 $X=221540 $Y=115060
X1049 1171 13 12 1598 79 1620 AO21X1 $T=237220 84100 0 180 $X=231400 $Y=78280
X1050 1161 13 12 1449 390 371 AO21X1 $T=237800 125860 0 180 $X=231980 $Y=120040
X1051 374 13 12 1604 33 1621 AO21X1 $T=234320 146740 1 0 $X=233720 $Y=140920
X1052 1162 13 12 1449 380 373 AO21X1 $T=236060 115420 0 0 $X=235460 $Y=115060
X1053 801 13 12 1622 1605 1288 AO21X1 $T=249400 146740 0 180 $X=243580 $Y=140920
X1054 1161 13 12 1450 1578 1623 AO21X1 $T=247080 125860 0 0 $X=246480 $Y=125500
X1055 379 13 12 1623 33 1624 AO21X1 $T=247660 115420 0 0 $X=247060 $Y=115060
X1056 631 13 12 1625 1626 1186 AO21X1 $T=256360 73660 1 180 $X=250540 $Y=73300
X1057 1162 13 12 1450 383 399 AO21X1 $T=253460 136300 1 0 $X=252860 $Y=130480
X1058 819 13 12 391 822 1344 AO21X1 $T=259840 52780 1 180 $X=254020 $Y=52420
X1059 820 13 12 398 823 1342 AO21X1 $T=264480 63220 0 180 $X=258660 $Y=57400
X1060 1181 13 12 615 808 387 AO21X1 $T=260420 31900 1 0 $X=259820 $Y=26080
X1061 1162 13 12 815 399 1386 AO21X1 $T=267380 125860 0 180 $X=261560 $Y=120040
X1062 634 13 12 1627 801 1628 AO21X1 $T=280140 84100 1 0 $X=279540 $Y=78280
X1063 1179 13 12 116 117 1313 AO21X1 $T=294640 178060 1 0 $X=294040 $Y=172240
X1064 115 13 12 870 1585 1629 AO21X1 $T=330020 167620 0 180 $X=324200 $Y=161800
X1065 1461 13 12 1629 108 1630 AO21X1 $T=332920 178060 0 0 $X=332320 $Y=177700
X1066 1210 13 12 882 1587 1631 AO21X1 $T=342780 157180 1 0 $X=342180 $Y=151360
X1067 892 13 12 1535 1211 1588 AO21X1 $T=352640 31900 0 180 $X=346820 $Y=26080
X1068 1462 13 12 1631 124 1632 AO21X1 $T=348000 157180 1 0 $X=347400 $Y=151360
X1069 893 13 12 1539 1212 1589 AO21X1 $T=357860 21460 1 180 $X=352040 $Y=21100
X1070 633 13 12 1599 124 1633 AO21X1 $T=366560 84100 1 180 $X=360740 $Y=83740
X1071 616 13 12 1634 1635 1236 AO21X1 $T=369460 84100 1 0 $X=368860 $Y=78280
X1072 1209 13 12 479 482 491 AO21X1 $T=381640 136300 1 0 $X=381040 $Y=130480
X1073 488 13 12 1636 108 1637 AO21X1 $T=383960 136300 0 0 $X=383360 $Y=135940
X1074 1201 13 12 1209 501 1316 AO21X1 $T=392660 115420 1 180 $X=386840 $Y=115060
X1075 1209 13 12 483 1592 1636 AO21X1 $T=390340 146740 0 0 $X=389740 $Y=146380
X1076 1209 13 12 1467 496 501 AO21X1 $T=392660 115420 0 0 $X=392060 $Y=115060
X1077 895 13 12 1209 496 1542 AO21X1 $T=393820 125860 1 0 $X=393220 $Y=120040
X1078 1210 13 12 1467 500 505 AO21X1 $T=397880 115420 0 0 $X=397280 $Y=115060
X1079 124 13 12 1638 1607 1304 AO21X1 $T=398460 167620 1 0 $X=397860 $Y=161800
X1080 504 13 12 499 491 1612 AO21X1 $T=402520 125860 0 0 $X=401920 $Y=125500
X1081 1238 13 12 1600 138 1639 AO21X1 $T=408900 94540 1 0 $X=408300 $Y=88720
X1082 1233 13 12 1640 1543 525 AO21X1 $T=415860 84100 0 0 $X=415260 $Y=83740
X1083 948 13 12 142 551 1320 AO21X1 $T=457620 178060 1 180 $X=451800 $Y=177700
X1084 142 13 12 166 169 542 AO21X1 $T=453560 188500 1 0 $X=452960 $Y=182680
X1085 988 13 12 142 170 173 AO21X1 $T=458780 188500 1 0 $X=458180 $Y=182680
X1086 144 13 12 1501 172 559 AO21X1 $T=460520 178060 1 0 $X=459920 $Y=172240
X1087 142 13 12 1501 170 551 AO21X1 $T=460520 178060 0 0 $X=459920 $Y=177700
X1088 1252 13 12 1548 993 1371 AO21X1 $T=484880 21460 1 180 $X=479060 $Y=21100
X1089 1253 13 12 1547 994 1377 AO21X1 $T=488360 31900 1 0 $X=487760 $Y=26080
X1090 1258 13 12 1602 186 1641 AO21X1 $T=502860 146740 1 0 $X=502260 $Y=140920
X1091 1263 13 12 1642 1569 194 AO21X1 $T=523160 157180 0 180 $X=517340 $Y=151360
X1092 47 43 13 12 42 XNOR2X1 $T=106140 188500 0 180 $X=99160 $Y=182680
X1093 420 49 13 12 1162 XNOR2X1 $T=190820 146740 1 180 $X=183840 $Y=146380
X1094 375 769 13 12 776 XNOR2X1 $T=233740 21460 1 180 $X=226760 $Y=21100
X1095 907 613 13 12 806 XNOR2X1 $T=276660 146740 1 180 $X=269680 $Y=146380
X1096 1231 116 13 12 1209 XNOR2X1 $T=366560 178060 0 180 $X=359580 $Y=172240
X1097 623 909 13 12 905 XNOR2X1 $T=375840 146740 1 180 $X=368860 $Y=146380
X1098 1248 1224 13 12 1222 XNOR2X1 $T=400200 31900 0 180 $X=393220 $Y=26080
X1099 1254 936 13 12 952 XNOR2X1 $T=458200 21460 1 180 $X=451220 $Y=21100
X1100 177 622 13 12 168 XNOR2X1 $T=480820 167620 1 180 $X=473840 $Y=167260
X1101 1272 1260 13 12 1261 XNOR2X1 $T=520260 31900 0 180 $X=513280 $Y=26080
X1102 1102 13 12 680 247 250 1125 OAI31XL $T=78880 115420 0 0 $X=78280 $Y=115060
X1103 628 13 12 686 1404 1615 706 OAI31XL $T=101500 115420 0 0 $X=100900 $Y=115060
X1104 1121 13 12 48 1333 261 1143 OAI31XL $T=115420 94540 0 0 $X=114820 $Y=94180
X1105 627 13 12 1124 1334 1616 730 OAI31XL $T=128180 104980 0 0 $X=127580 $Y=104620
X1106 33 13 12 283 281 1617 66 OAI31XL $T=149060 188500 1 0 $X=148460 $Y=182680
X1107 312 13 12 310 1643 1618 440 OAI31XL $T=167040 146740 1 180 $X=161800 $Y=146380
X1108 754 13 12 1158 338 1619 775 OAI31XL $T=203580 94540 0 0 $X=202980 $Y=94180
X1109 1171 13 12 1168 1343 1620 802 OAI31XL $T=226780 84100 1 0 $X=226180 $Y=78280
X1110 362 13 12 378 1644 1621 1197 OAI31XL $T=239540 146740 1 0 $X=238940 $Y=140920
X1111 801 13 12 390 400 1624 1287 OAI31XL $T=255780 125860 1 0 $X=255180 $Y=120040
X1112 634 13 12 1185 417 1628 866 OAI31XL $T=291160 84100 1 0 $X=290560 $Y=78280
X1113 837 13 12 834 429 1193 1349 OAI31XL $T=309720 42340 1 180 $X=304480 $Y=41980
X1114 836 13 12 833 435 1192 1348 OAI31XL $T=314360 42340 1 180 $X=309120 $Y=41980
X1115 427 13 12 123 1645 124 1646 OAI31XL $T=310300 188500 1 0 $X=309700 $Y=182680
X1116 124 13 12 125 1314 1646 472 OAI31XL $T=316100 178060 1 180 $X=310860 $Y=177700
X1117 124 13 12 456 453 1630 129 OAI31XL $T=338140 178060 0 0 $X=337540 $Y=177700
X1118 1218 13 12 1216 1588 1214 1352 OAI31XL $T=353220 42340 0 180 $X=347980 $Y=36520
X1119 108 13 12 1537 1565 1632 1297 OAI31XL $T=350900 157180 0 0 $X=350300 $Y=156820
X1120 1219 13 12 1217 1589 1215 1353 OAI31XL $T=359600 42340 0 180 $X=354360 $Y=36520
X1121 633 13 12 1221 1356 1633 911 OAI31XL $T=368300 84100 0 180 $X=363060 $Y=78280
X1122 486 13 12 491 1647 108 1648 OAI31XL $T=382800 115420 1 0 $X=382200 $Y=109600
X1123 124 13 12 482 1567 1637 1305 OAI31XL $T=385120 146740 1 0 $X=384520 $Y=140920
X1124 108 13 12 490 1317 1648 497 OAI31XL $T=389180 125860 1 0 $X=388580 $Y=120040
X1125 1238 13 12 1235 508 1639 928 OAI31XL $T=407740 94540 0 180 $X=402500 $Y=88720
X1126 137 13 12 160 1321 1649 158 OAI31XL $T=443700 188500 0 180 $X=438460 $Y=182680
X1127 540 13 12 542 1650 137 1649 OAI31XL $T=444280 178060 0 180 $X=439040 $Y=172240
X1128 1258 13 12 1030 1379 1641 1056 OAI31XL $T=494740 146740 1 0 $X=494140 $Y=140920
X1129 1099 1105 13 12 245 1107 1402 AOI31XL $T=78300 73660 0 0 $X=77700 $Y=73300
X1130 1106 1100 13 12 251 1108 253 AOI31XL $T=90480 73660 0 0 $X=89880 $Y=73300
X1131 304 311 13 12 1427 33 1425 AOI31XL $T=158340 157180 1 0 $X=157740 $Y=151360
X1132 77 1151 13 12 326 1527 344 AOI31XL $T=190240 84100 1 0 $X=189640 $Y=78280
X1133 372 361 13 12 1439 801 1441 AOI31XL $T=233740 136300 1 180 $X=228500 $Y=135940
X1134 79 778 13 12 370 1625 401 AOI31XL $T=252300 73660 1 0 $X=251700 $Y=67840
X1135 122 426 13 12 120 108 1459 AOI31XL $T=304500 188500 1 0 $X=303900 $Y=182680
X1136 852 1188 13 12 433 1533 446 AOI31XL $T=305660 84100 1 0 $X=305060 $Y=78280
X1137 124 1207 13 12 459 1634 475 AOI31XL $T=357280 84100 1 0 $X=356680 $Y=78280
X1138 492 485 13 12 1479 124 1476 AOI31XL $T=387440 104980 0 0 $X=386840 $Y=104620
X1139 138 922 13 12 517 1640 519 AOI31XL $T=414700 84100 1 0 $X=414100 $Y=78280
X1140 543 539 13 12 1497 138 1487 AOI31XL $T=450080 167620 1 180 $X=444840 $Y=167260
X1141 186 1035 13 12 575 578 583 AOI31XL $T=505180 125860 1 0 $X=504580 $Y=120040
X1142 30 53 13 12 1608 296 1553 AOI211XL $T=149640 178060 0 180 $X=144980 $Y=172240
X1143 1127 53 13 12 1392 291 1555 AOI211XL $T=150220 157180 1 180 $X=145560 $Y=156820
X1144 1166 1162 13 12 1394 373 1559 AOI211XL $T=240120 125860 1 180 $X=235460 $Y=125500
X1145 816 1162 13 12 1609 380 1561 AOI211XL $T=247080 104980 1 180 $X=242420 $Y=104620
X1146 899 1210 13 12 1610 487 495 AOI211XL $T=392660 136300 0 180 $X=388000 $Y=130480
X1147 1199 1210 13 12 1611 490 502 AOI211XL $T=403100 125860 0 180 $X=398440 $Y=120040
X1148 986 144 13 12 1613 160 552 AOI211XL $T=460520 178060 0 180 $X=455860 $Y=172240
X1149 31 13 12 655 236 238 1399 654 AOI32XL $T=69020 52780 1 180 $X=63200 $Y=52420
X1150 727 13 12 1142 302 318 308 729 AOI32XL $T=165300 94540 1 180 $X=159480 $Y=94180
X1151 1242 13 12 1244 536 555 547 151 AOI32XL $T=451240 104980 1 0 $X=450640 $Y=99160
X1152 671 13 12 711 1570 231 ACHCONX2 $T=48140 157180 0 0 $X=47560 $Y=156820
X1153 28 13 12 30 242 36 ACHCONX2 $T=50460 188500 1 0 $X=49880 $Y=182680
X1154 26 13 12 29 34 248 ACHCONX2 $T=52200 178060 0 0 $X=51620 $Y=177700
X1155 711 13 12 670 1571 243 ACHCONX2 $T=55100 167620 1 0 $X=54520 $Y=161800
X1156 1126 13 12 683 1651 1570 ACHCONX2 $T=77140 157180 1 0 $X=76560 $Y=151360
X1157 1126 13 12 684 1652 1571 ACHCONX2 $T=77140 157180 0 0 $X=76560 $Y=156820
X1158 709 13 12 1132 1572 1651 ACHCONX2 $T=108460 136300 1 0 $X=107880 $Y=130480
X1159 1132 13 12 708 297 1652 ACHCONX2 $T=108460 136300 0 0 $X=107880 $Y=135940
X1160 732 13 12 715 1573 298 ACHCONX2 $T=128760 125860 0 0 $X=128180 $Y=125500
X1161 731 13 12 715 322 1572 ACHCONX2 $T=130500 125860 1 0 $X=129920 $Y=120040
X1162 731 13 12 53 1643 1427 ACHCONX2 $T=150220 146740 1 0 $X=149640 $Y=140920
X1163 68 13 12 49 284 1574 ACHCONX2 $T=158920 178060 0 0 $X=158340 $Y=177700
X1164 607 13 12 1162 1578 322 ACHCONX2 $T=165880 125860 1 0 $X=165300 $Y=120040
X1165 607 13 12 1161 383 1573 ACHCONX2 $T=165880 125860 0 0 $X=165300 $Y=125500
X1166 762 13 12 774 78 342 ACHCONX2 $T=167040 157180 1 0 $X=166460 $Y=151360
X1167 763 13 12 774 1574 333 ACHCONX2 $T=167040 157180 0 0 $X=166460 $Y=156820
X1168 765 13 12 1166 1577 358 ACHCONX2 $T=198360 104980 0 0 $X=197780 $Y=104620
X1169 764 13 12 1166 353 352 ACHCONX2 $T=198360 125860 1 0 $X=197780 $Y=120040
X1170 1163 13 12 766 333 1577 ACHCONX2 $T=227360 136300 1 180 $X=197780 $Y=135940
X1171 1164 13 12 766 341 354 ACHCONX2 $T=198360 146740 0 0 $X=197780 $Y=146380
X1172 773 13 12 1162 1644 1439 ACHCONX2 $T=210540 157180 1 0 $X=209960 $Y=151360
X1173 1161 13 12 806 1622 1578 ACHCONX2 $T=224460 136300 1 0 $X=223880 $Y=130480
X1174 817 13 12 797 351 404 ACHCONX2 $T=259260 94540 1 180 $X=229680 $Y=94180
X1175 803 13 12 1180 1582 411 ACHCONX2 $T=246500 167620 1 0 $X=245920 $Y=161800
X1176 793 13 12 96 410 409 ACHCONX2 $T=246500 178060 0 0 $X=245920 $Y=177700
X1177 799 13 12 104 1579 106 ACHCONX2 $T=247080 188500 1 0 $X=246500 $Y=182680
X1178 804 13 12 1180 1581 412 ACHCONX2 $T=254620 157180 0 0 $X=254040 $Y=156820
X1179 818 13 12 797 357 414 ACHCONX2 $T=256940 104980 0 0 $X=256360 $Y=104620
X1180 828 13 12 816 403 423 ACHCONX2 $T=256940 115420 1 0 $X=256360 $Y=109600
X1181 828 13 12 815 414 1580 ACHCONX2 $T=256940 115420 0 0 $X=256360 $Y=115060
X1182 814 13 12 812 1580 1532 ACHCONX2 $T=256940 136300 0 0 $X=256360 $Y=135940
X1183 97 13 12 793 412 1579 ACHCONX2 $T=256940 178060 1 0 $X=256360 $Y=172240
X1184 813 13 12 812 422 1531 ACHCONX2 $T=288260 146740 1 0 $X=287680 $Y=140920
X1185 848 13 12 115 1645 120 ACHCONX2 $T=288260 167620 0 0 $X=287680 $Y=167260
X1186 848 13 12 842 1564 1581 ACHCONX2 $T=295800 167620 1 0 $X=295220 $Y=161800
X1187 845 13 12 1202 1583 449 ACHCONX2 $T=298700 104980 0 0 $X=298120 $Y=104620
X1188 868 13 12 860 1585 1583 ACHCONX2 $T=303920 125860 0 0 $X=303340 $Y=125500
X1189 843 13 12 848 1587 1582 ACHCONX2 $T=305080 157180 1 0 $X=304500 $Y=151360
X1190 1198 13 12 854 450 1590 ACHCONX2 $T=313780 94540 1 0 $X=313200 $Y=88720
X1191 846 13 12 1202 1584 450 ACHCONX2 $T=313780 115420 1 0 $X=313200 $Y=109600
X1192 860 13 12 867 1586 1584 ACHCONX2 $T=313780 125860 1 0 $X=313200 $Y=120040
X1193 854 13 12 1199 448 454 ACHCONX2 $T=314360 94540 0 0 $X=313780 $Y=94180
X1194 128 13 12 115 1653 1629 ACHCONX2 $T=343940 188500 0 180 $X=314360 $Y=182680
X1195 885 13 12 1210 1654 1631 ACHCONX2 $T=338140 146740 1 0 $X=337560 $Y=140920
X1196 895 13 12 902 454 1591 ACHCONX2 $T=341620 104980 1 0 $X=341040 $Y=99160
X1197 902 13 12 896 1590 471 ACHCONX2 $T=344520 94540 1 0 $X=343940 $Y=88720
X1198 889 13 12 899 470 1540 ACHCONX2 $T=346260 125860 1 0 $X=345680 $Y=120040
X1199 860 13 12 1210 1647 1479 ACHCONX2 $T=346840 115420 1 0 $X=346260 $Y=109600
X1200 899 13 12 888 1591 1538 ACHCONX2 $T=346840 125860 0 0 $X=346260 $Y=125500
X1201 916 13 12 1209 1638 1592 ACHCONX2 $T=378160 167620 0 0 $X=377580 $Y=167260
X1202 939 13 12 148 153 524 ACHCONX2 $T=399040 178060 1 0 $X=398460 $Y=172240
X1203 940 13 12 148 156 527 ACHCONX2 $T=407160 167620 0 0 $X=406580 $Y=167260
X1204 943 13 12 949 1593 1655 ACHCONX2 $T=408900 136300 1 0 $X=408320 $Y=130480
X1205 945 13 12 929 527 1593 ACHCONX2 $T=410060 146740 1 0 $X=409480 $Y=140920
X1206 929 13 12 946 523 538 ACHCONX2 $T=412960 136300 0 0 $X=412380 $Y=135940
X1207 942 13 12 949 537 1656 ACHCONX2 $T=428040 125860 1 0 $X=427460 $Y=120040
X1208 945 13 12 144 1650 1497 ACHCONX2 $T=428620 167620 1 0 $X=428040 $Y=161800
X1209 985 13 12 983 1656 1594 ACHCONX2 $T=465740 125860 1 180 $X=436160 $Y=125500
X1210 985 13 12 982 1655 1595 ACHCONX2 $T=468060 136300 1 0 $X=467480 $Y=130480
X1211 1017 13 12 989 1594 1545 ACHCONX2 $T=468060 146740 0 0 $X=467480 $Y=146380
X1212 1018 13 12 989 1595 1546 ACHCONX2 $T=468060 157180 1 0 $X=467480 $Y=151360
X1213 1026 13 12 179 581 187 ACHCONX2 $T=479080 188500 1 0 $X=478500 $Y=182680
X1214 180 13 12 181 587 188 ACHCONX2 $T=489520 178060 1 0 $X=488940 $Y=172240
X1215 185 13 12 181 197 582 ACHCONX2 $T=502280 178060 0 0 $X=501700 $Y=177700
X1216 1063 13 12 192 198 587 ACHCONX2 $T=505760 167620 0 0 $X=505180 $Y=167260
X1217 1313 13 12 121 1315 108 1460 AND4XL $T=305660 178060 0 0 $X=305060 $Y=177700
X1218 1316 13 12 489 1319 124 1477 AND4XL $T=382220 125860 1 0 $X=381620 $Y=120040
X1219 1601 13 12 1242 1244 1239 1485 AND4XL $T=433260 94540 0 0 $X=432660 $Y=94180
X1220 1320 13 12 541 1323 138 1488 AND4XL $T=447760 178060 1 180 $X=441940 $Y=177700
X1221 558 13 12 1249 1020 1255 1508 AND4XL $T=480240 115420 1 0 $X=479640 $Y=109600
X1222 1657 13 12 1266 1268 1065 1642 AND4XL $T=528960 125860 1 180 $X=523140 $Y=125500
X1223 1658 13 12 1082 1068 1085 1657 AND4XL $T=533600 94540 1 180 $X=527780 $Y=94180
X1224 1659 13 12 1076 1079 1091 1658 AND4XL $T=529540 73660 1 0 $X=528940 $Y=67840
X1225 1073 13 12 1071 1088 1270 1659 AND4XL $T=536500 52780 1 180 $X=530680 $Y=52420
X1226 1366 1244 13 12 975 972 1489 OR4XL $T=448920 94540 0 180 $X=443100 $Y=88720
X1227 1660 1065 13 12 1268 1266 1568 OR4XL $T=522580 125860 1 180 $X=516760 $Y=125500
X1228 1661 1091 13 12 1079 1076 1662 OR4XL $T=529540 73660 0 180 $X=523720 $Y=67840
X1229 1662 1082 13 12 1085 1068 1660 OR4XL $T=531280 104980 0 180 $X=525460 $Y=99160
X1230 1071 1073 13 12 1270 1088 1661 OR4XL $T=539400 52780 0 180 $X=533580 $Y=46960
X1231 40 13 12 1596 249 685 630 AO22X1 $T=91640 115420 1 180 $X=85240 $Y=115060
X1232 1157 13 12 1528 1597 72 1172 AO22X1 $T=198360 94540 1 0 $X=197760 $Y=88720
X1233 1167 13 12 1626 1598 93 1183 AO22X1 $T=243020 84100 0 180 $X=236620 $Y=78280
X1234 1184 13 12 1533 1627 33 636 AO22X1 $T=278400 84100 0 180 $X=272000 $Y=78280
X1235 1220 13 12 1635 1599 108 477 AO22X1 $T=368300 84100 0 0 $X=367700 $Y=83740
X1236 1234 13 12 1543 1600 137 1241 AO22X1 $T=405420 84100 0 0 $X=404820 $Y=83740
X1237 1029 13 12 574 1602 183 1265 AO22X1 $T=504600 136300 0 0 $X=504000 $Y=135940
X1238 419 851 13 12 1187 825 416 AND4X1 $T=294060 73660 1 180 $X=288240 $Y=73300
X1239 1534 1188 13 12 1185 852 1627 AND4X1 $T=303340 84100 0 180 $X=297520 $Y=78280
X1240 564 1057 13 12 1041 1044 569 AND4X1 $T=499960 52780 0 0 $X=499360 $Y=52420
X1241 1418 1141 13 12 726 1136 1557 OR4X1 $T=146160 104980 1 0 $X=145560 $Y=99160
X1242 1338 727 13 12 1142 721 307 OR4X1 $T=147320 94540 1 0 $X=146720 $Y=88720
X1243 1518 1041 13 12 1057 1044 1382 OR4X1 $T=519100 52780 1 180 $X=513280 $Y=52420
X1244 734 729 13 12 735 64 736 1156 733 OAI222XL $T=174000 42340 0 180 $X=167020 $Y=36520
X1245 1124 1411 13 12 264 705 273 OA22X1 $T=118320 115420 1 0 $X=117720 $Y=109600
X1246 311 1414 13 12 53 NAND2BX1 $T=156600 157180 0 0 $X=156000 $Y=156820
X1247 1153 1339 13 12 302 NAND2BX1 $T=157760 84100 0 0 $X=157160 $Y=83740
X1248 361 1435 13 12 1162 NAND2BX1 $T=222720 136300 0 180 $X=218640 $Y=130480
X1249 432 1534 13 12 801 NAND2BX1 $T=306820 73660 0 180 $X=302740 $Y=67840
X1250 127 1461 13 12 1653 NAND2BX1 $T=327120 178060 0 0 $X=326520 $Y=177700
X1251 1566 1462 13 12 1654 NAND2BX1 $T=348000 146740 0 0 $X=347400 $Y=146380
X1252 481 1469 13 12 1210 NAND2BX1 $T=379320 146740 1 0 $X=378720 $Y=140920
X1253 535 1601 13 12 151 NAND2BX1 $T=440220 94540 0 0 $X=439620 $Y=94180
X1254 33 1651 13 12 1652 1275 MX2X1 $T=113100 146740 0 0 $X=112500 $Y=146380
X1255 33 1531 13 12 1532 1291 MX2X1 $T=297540 125860 1 180 $X=291720 $Y=125500
X1256 108 1538 13 12 1540 1300 MX2X1 $T=373520 136300 0 180 $X=367700 $Y=130480
X1257 137 1656 13 12 1655 1309 MX2X1 $T=460520 136300 0 180 $X=454700 $Y=130480
X1258 137 1545 13 12 1546 1311 MX2X1 $T=475020 157180 0 0 $X=474420 $Y=156820
X1259 1561 13 12 1623 816 1162 AOI2BB1X1 $T=247660 115420 1 180 $X=242420 $Y=115060
X1260 495 13 12 1636 899 1210 AOI2BB1X1 $T=389180 136300 0 0 $X=388580 $Y=135940
X1261 1663 13 12 542 1614 172 AOI2BB1X1 $T=468060 178060 0 0 $X=467460 $Y=177700
X1262 1138 13 12 1411 701 260 OAI2BB1X1 $T=122960 104980 0 180 $X=118300 $Y=99160
X1263 452 13 12 1586 870 116 OAI2BB1X1 $T=342200 157180 1 180 $X=337540 $Y=156820
X1264 1404 40 249 13 12 NOR2XL $T=85840 115420 1 180 $X=82920 $Y=115060
X1265 1343 93 1626 13 12 NOR2XL $T=241280 73660 0 0 $X=240680 $Y=73300
X1266 1356 108 1635 13 12 NOR2XL $T=370620 73660 0 0 $X=370020 $Y=73300
X1267 1663 174 13 12 INVXL $T=468060 188500 1 0 $X=467460 $Y=182680
X1268 33 13 12 1556 1424 1526 292 NOR4BBX1 $T=150220 157180 1 0 $X=149620 $Y=151360
X1269 801 13 12 1560 1440 1529 374 NOR4BBX1 $T=223300 146740 1 0 $X=222700 $Y=140920
X1270 1530 13 12 93 1625 AND2X1 $T=245920 73660 0 0 $X=245320 $Y=73300
X1271 1347 13 12 432 438 AND2X1 $T=311460 73660 1 0 $X=310860 $Y=67840
X1272 1536 13 12 108 1634 AND2X1 $T=352640 84100 1 0 $X=352040 $Y=78280
X1273 1544 13 12 137 1640 AND2X1 $T=421080 84100 0 0 $X=420480 $Y=83740
.ends MASCO__P1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ADDFXL                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ADDFXL CO VDD VSS B A CI S
** N=19 EP=7 FDC=28
M0 CO 9 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=710 $Y=1290 $dt=0
M1 VSS A 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2690 $Y=1360 $dt=0
M2 10 B VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3530 $Y=1320 $dt=0
M3 9 CI 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4370 $Y=1320 $dt=0
M4 11 B 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=6570 $Y=800 $dt=0
M5 VSS A 11 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7010 $Y=800 $dt=0
M6 12 CI VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7850 $Y=800 $dt=0
M7 VSS B 12 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=8690 $Y=800 $dt=0
M8 12 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=9770 $Y=800 $dt=0
M9 8 9 12 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=10610 $Y=800 $dt=0
M10 13 CI 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=12230 $Y=800 $dt=0
M11 14 B 13 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=12670 $Y=800 $dt=0
M12 VSS A 14 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=13110 $Y=800 $dt=0
M13 S 8 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=13950 $Y=800 $dt=0
M14 CO 9 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=710 $Y=3450 $dt=1
M15 VDD A 15 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2690 $Y=2800 $dt=1
M16 15 B VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3530 $Y=3080 $dt=1
M17 9 CI 15 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4370 $Y=3080 $dt=1
M18 16 B 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=6020 $Y=3340 $dt=1
M19 VDD A 16 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=6520 $Y=3340 $dt=1
M20 17 CI VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7360 $Y=3040 $dt=1
M21 VDD B 17 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=8200 $Y=3040 $dt=1
M22 17 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=9040 $Y=3520 $dt=1
M23 8 9 17 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=10120 $Y=3520 $dt=1
M24 18 CI 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=11740 $Y=3700 $dt=1
M25 19 B 18 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=12180 $Y=3700 $dt=1
M26 VDD A 19 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=12620 $Y=3700 $dt=1
M27 S 8 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=13700 $Y=3700 $dt=1
.ends ADDFXL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MXI3X1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MXI3X1 S0 A VDD VSS B S1 C Y
** N=21 EP=8 FDC=24
M0 VSS S0 13 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1030 $Y=1240 $dt=0
M1 14 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1870 $Y=1240 $dt=0
M2 12 13 14 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2310 $Y=1240 $dt=0
M3 15 S0 12 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3150 $Y=1240 $dt=0
M4 VSS B 15 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4150 $Y=1240 $dt=0
M5 16 12 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4990 $Y=1240 $dt=0
M6 9 11 16 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5430 $Y=1240 $dt=0
M7 17 S1 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=6910 $Y=1240 $dt=0
M8 VSS 10 17 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7630 $Y=1240 $dt=0
M9 11 S1 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=8470 $Y=1240 $dt=0
M10 VSS C 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=10090 $Y=1080 $dt=0
M11 Y 9 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=10930 $Y=980 $dt=0
M12 VDD S0 13 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1190 $Y=3360 $dt=1
M13 18 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2030 $Y=3360 $dt=1
M14 12 S0 18 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2830 $Y=3360 $dt=1
M15 19 13 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3670 $Y=3360 $dt=1
M16 VDD B 19 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4150 $Y=3360 $dt=1
M17 20 12 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5110 $Y=3360 $dt=1
M18 9 S1 20 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5550 $Y=3360 $dt=1
M19 21 11 9 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=6470 $Y=3360 $dt=1
M20 VDD 10 21 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=6990 $Y=3360 $dt=1
M21 11 S1 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=8070 $Y=3360 $dt=1
M22 VDD C 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=9850 $Y=2680 $dt=1
M23 Y 9 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=10930 $Y=2680 $dt=1
.ends MXI3X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: SDFFRX1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt SDFFRX1 QN VDD VSS Q CK RN D SI SE
** N=28 EP=9 FDC=40
M0 VSS 17 QN VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=980 $dt=0
M1 17 15 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1550 $Y=1360 $dt=0
M2 VSS 15 Q VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=3170 $Y=980 $dt=0
M3 11 CK VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4130 $Y=1360 $dt=0
M4 18 16 15 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=6130 $Y=1240 $dt=0
M5 VSS RN 18 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=6570 $Y=1240 $dt=0
M6 19 15 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=7650 $Y=1240 $dt=0
M7 16 11 19 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=8370 $Y=1240 $dt=0
M8 13 12 16 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=9970 $Y=1240 $dt=0
M9 VSS 14 13 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=11010 $Y=1240 $dt=0
M10 20 RN VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=12210 $Y=1240 $dt=0
M11 21 13 20 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=12650 $Y=1240 $dt=0
M12 14 12 21 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=13370 $Y=1240 $dt=0
M13 22 11 14 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=14210 $Y=1240 $dt=0
M14 VSS 11 12 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=15970 $Y=800 $dt=0
M15 23 D VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=17090 $Y=800 $dt=0
M16 22 10 23 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=17970 $Y=800 $dt=0
M17 24 SE 22 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=18810 $Y=800 $dt=0
M18 VSS SI 24 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=19250 $Y=800 $dt=0
M19 10 SE VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=20090 $Y=800 $dt=0
M20 VDD 17 QN VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=710 $Y=2680 $dt=1
M21 17 15 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1550 $Y=2680 $dt=1
M22 VDD 15 Q VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=3170 $Y=3120 $dt=1
M23 11 CK VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4130 $Y=3120 $dt=1
M24 15 16 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=5730 $Y=3020 $dt=1
M25 VDD RN 15 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=6570 $Y=3020 $dt=1
M26 25 15 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=7650 $Y=3020 $dt=1
M27 16 12 25 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=8530 $Y=3020 $dt=1
M28 13 11 16 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=9530 $Y=3020 $dt=1
M29 VDD 14 13 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=10570 $Y=3020 $dt=1
M30 26 RN VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=11650 $Y=3020 $dt=1
M31 VDD 13 26 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=12490 $Y=3020 $dt=1
M32 14 11 26 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=13990 $Y=2680 $dt=1
M33 22 12 14 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=14830 $Y=2680 $dt=1
M34 VDD 11 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=16450 $Y=3180 $dt=1
M35 27 D VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=17290 $Y=3180 $dt=1
M36 22 SE 27 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=17730 $Y=3180 $dt=1
M37 28 10 22 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=18570 $Y=3180 $dt=1
M38 VDD SI 28 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=19050 $Y=3180 $dt=1
M39 10 SE VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=19890 $Y=3180 $dt=1
.ends SDFFRX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR3XL                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR3XL A B VDD VSS C Y
** N=13 EP=6 FDC=22
M0 VSS A 10 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=970 $Y=800 $dt=0
M1 11 B VSS VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=2050 $Y=800 $dt=0
M2 9 10 VSS VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=4410 $Y=800 $dt=0
M3 12 11 9 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=5490 $Y=800 $dt=0
M4 10 B 12 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=7090 $Y=800 $dt=0
M5 13 11 10 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=8170 $Y=800 $dt=0
M6 9 B 13 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=9500 $Y=800 $dt=0
M7 7 C 12 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=12120 $Y=800 $dt=0
M8 13 8 7 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=13200 $Y=800 $dt=0
M9 VSS C 8 VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=15060 $Y=800 $dt=0
M10 Y 7 VSS VSS nmos1v L=1e-07 W=3.2e-07 fw=3.2e-07 simw=3.2e-07 $X=16140 $Y=800 $dt=0
M11 VDD A 10 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=970 $Y=3380 $dt=1
M12 11 B VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=2050 $Y=3380 $dt=1
M13 9 10 VDD VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=4410 $Y=3380 $dt=1
M14 12 B 9 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=5490 $Y=3380 $dt=1
M15 10 11 12 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=6650 $Y=3340 $dt=1
M16 13 B 10 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=8150 $Y=2940 $dt=1
M17 9 11 13 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=9230 $Y=3340 $dt=1
M18 7 8 12 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=12120 $Y=3380 $dt=1
M19 13 C 7 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=13200 $Y=3380 $dt=1
M20 VDD C 8 VDD pmos1v L=1e-07 W=5.2e-07 fw=5.2e-13 simw=5.2e-07 $X=15060 $Y=3380 $dt=1
M21 Y 7 VDD VDD pmos1v L=1e-07 W=3.4e-07 fw=3.4e-13 simw=3.4e-07 $X=16140 $Y=3740 $dt=1
.ends XOR3XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: CLKXOR2X1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt CLKXOR2X1 Y VDD VSS A B
** N=10 EP=5 FDC=12
M0 VSS 8 Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=980 $dt=0
M1 6 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1830 $Y=1080 $dt=0
M2 8 7 6 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3110 $Y=1080 $dt=0
M3 9 B 8 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3950 $Y=1080 $dt=0
M4 VSS 6 9 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4390 $Y=1080 $dt=0
M5 7 B VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5230 $Y=1080 $dt=0
M6 VDD 8 Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=780 $Y=3120 $dt=1
M7 6 A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1860 $Y=3240 $dt=1
M8 8 B 6 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2700 $Y=3240 $dt=1
M9 10 7 8 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3540 $Y=3240 $dt=1
M10 VDD 6 10 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4150 $Y=3240 $dt=1
M11 7 B VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4990 $Y=3240 $dt=1
.ends CLKXOR2X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OAI21X1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OAI21X1 A0 A1 VDD VSS B0 Y
** N=8 EP=6 FDC=6
M0 VSS A0 7 VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=890 $Y=800 $dt=0
M1 7 A1 VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1730 $Y=800 $dt=0
M2 Y B0 7 VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=2570 $Y=800 $dt=0
M3 8 A0 VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1290 $Y=3120 $dt=1
M4 Y A1 8 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1730 $Y=3120 $dt=1
M5 VDD B0 Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=2570 $Y=3120 $dt=1
.ends OAI21X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NOR3BX1                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NOR3BX1 C Y B VDD VSS AN
** N=9 EP=6 FDC=8
M0 VSS C Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=800 $dt=0
M1 Y B VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1550 $Y=800 $dt=0
M2 VSS 7 Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=2390 $Y=800 $dt=0
M3 7 AN VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3230 $Y=800 $dt=0
M4 8 C Y VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1190 $Y=3120 $dt=1
M5 9 B 8 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1630 $Y=3120 $dt=1
M6 VDD 7 9 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=2270 $Y=3120 $dt=1
M7 7 AN VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3230 $Y=3120 $dt=1
.ends NOR3BX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NOR3X1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NOR3X1 A VDD VSS Y B C
** N=8 EP=6 FDC=6
M0 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=710 $Y=800 $dt=0
M1 VSS B Y VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=1550 $Y=800 $dt=0
M2 Y C VSS VSS nmos1v L=1e-07 W=4.3e-07 fw=4.3e-07 simw=4.3e-07 $X=2390 $Y=800 $dt=0
M3 7 A VDD VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=780 $Y=2900 $dt=1
M4 8 B 7 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=1420 $Y=2900 $dt=1
M5 Y C 8 VDD pmos1v L=1e-07 W=6.5e-07 fw=6.5e-13 simw=6.5e-07 $X=2060 $Y=2900 $dt=1
.ends NOR3X1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__P2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__P2 6 10 11 22 23 24 25 26 27 28
+ 29 30 31 32 33 34 35 36 37 38
+ 39 40 41 42 43 44 45 46 47 49
+ 50 51 52 54 55 56 57 58 59 60
+ 61 62 65 66 67 68 69 70 71 72
+ 73 74 75 76 77 78 80 82 83 84
+ 85 86 87 88 89 90 91 92 93 94
+ 95 96 97 98 99 100 101 102 103 104
+ 105 106 107 108 109 110 111 112 113 114
+ 115 116 117 118 119 120 121 122 123 124
+ 125 126 127 128 129 130 131 132 133 134
+ 135 136 137 138 139 140 141 142 143 144
+ 145 146 147 148 149 150 151 152 153 154
+ 155 156 157 158 159 160 161 162 163 164
+ 165 166 167 168 169 170 171 172 173 174
+ 175 176 178 179 180 181 182 183 184 185
+ 186 187 188 190 192 193 194 195 196 197
+ 198 199 200 201 202 203 204 205 206 207
+ 208 209 210 211 212 213 216 217 218 219
+ 220 221 222 224 225 226 227 228 229 231
+ 232 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252
+ 253 254 255 257 258 259 261 262 263 264
+ 265 267 268 269 270 271 272 273 274 276
+ 277 278 279 280 281 282 283 284 285 286
+ 287 288 289 291 292 293 294 295 297 298
+ 299 301 302 304 305 307 308 309 310 311
+ 313 314 315 316
** N=1832 EP=274 FDC=22396
X0 330 11 10 6 CLKBUFX2 $T=35380 365980 1 0 $X=34780 $Y=360160
X1 331 11 10 22 CLKBUFX2 $T=38860 365980 1 0 $X=38260 $Y=360160
X2 332 11 10 40 CLKBUFX2 $T=66120 355540 0 0 $X=65520 $Y=355180
X3 124 11 10 102 CLKINVX2 $T=372360 376420 1 0 $X=371760 $Y=370600
X4 124 11 10 221 CLKINVX2 $T=397880 376420 1 0 $X=397280 $Y=370600
X5 333 334 11 10 CLKINVX1 $T=60900 240700 1 180 $X=58560 $Y=240340
X6 335 336 11 10 CLKINVX1 $T=63220 230260 1 180 $X=60880 $Y=229900
X7 337 338 11 10 CLKINVX1 $T=71920 345100 0 0 $X=71320 $Y=344740
X8 339 340 11 10 CLKINVX1 $T=75400 188500 1 180 $X=73060 $Y=188140
X9 341 342 11 10 CLKINVX1 $T=75980 251140 0 0 $X=75380 $Y=250780
X10 46 49 11 10 CLKINVX1 $T=76560 188500 0 0 $X=75960 $Y=188140
X11 343 344 11 10 CLKINVX1 $T=78300 334660 0 180 $X=75960 $Y=328840
X12 345 346 11 10 CLKINVX1 $T=77720 272020 1 0 $X=77120 $Y=266200
X13 347 348 11 10 CLKINVX1 $T=84680 334660 0 180 $X=82340 $Y=328840
X14 349 350 11 10 CLKINVX1 $T=87000 292900 0 0 $X=86400 $Y=292540
X15 351 352 11 10 CLKINVX1 $T=91060 209380 1 180 $X=88720 $Y=209020
X16 353 354 11 10 CLKINVX1 $T=93960 209380 1 0 $X=93360 $Y=203560
X17 355 356 11 10 CLKINVX1 $T=98020 209380 1 180 $X=95680 $Y=209020
X18 357 358 11 10 CLKINVX1 $T=97440 219820 1 0 $X=96840 $Y=214000
X19 359 360 11 10 CLKINVX1 $T=97440 292900 0 0 $X=96840 $Y=292540
X20 361 362 11 10 CLKINVX1 $T=100920 219820 0 180 $X=98580 $Y=214000
X21 363 364 11 10 CLKINVX1 $T=99180 292900 0 0 $X=98580 $Y=292540
X22 365 366 11 10 CLKINVX1 $T=99760 334660 1 0 $X=99160 $Y=328840
X23 367 368 11 10 CLKINVX1 $T=103240 272020 0 180 $X=100900 $Y=266200
X24 369 370 11 10 CLKINVX1 $T=103820 324220 0 0 $X=103220 $Y=323860
X25 371 372 11 10 CLKINVX1 $T=108460 209380 1 0 $X=107860 $Y=203560
X26 373 374 11 10 CLKINVX1 $T=113100 292900 0 180 $X=110760 $Y=287080
X27 375 376 11 10 CLKINVX1 $T=116580 209380 1 0 $X=115980 $Y=203560
X28 377 378 11 10 CLKINVX1 $T=118320 209380 1 0 $X=117720 $Y=203560
X29 379 78 11 10 CLKINVX1 $T=125860 198940 1 180 $X=123520 $Y=198580
X30 380 381 11 10 CLKINVX1 $T=125860 292900 1 0 $X=125260 $Y=287080
X31 382 383 11 10 CLKINVX1 $T=133400 313780 1 180 $X=131060 $Y=313420
X32 384 385 11 10 CLKINVX1 $T=133980 209380 1 0 $X=133380 $Y=203560
X33 386 387 11 10 CLKINVX1 $T=134560 292900 0 0 $X=133960 $Y=292540
X34 388 389 11 10 CLKINVX1 $T=135720 219820 1 0 $X=135120 $Y=214000
X35 390 391 11 10 CLKINVX1 $T=137460 230260 0 0 $X=136860 $Y=229900
X36 392 393 11 10 CLKINVX1 $T=139200 324220 0 180 $X=136860 $Y=318400
X37 394 395 11 10 CLKINVX1 $T=140940 230260 1 180 $X=138600 $Y=229900
X38 396 397 11 10 CLKINVX1 $T=145580 219820 1 0 $X=144980 $Y=214000
X39 398 399 11 10 CLKINVX1 $T=151960 230260 0 180 $X=149620 $Y=224440
X40 400 401 11 10 CLKINVX1 $T=152540 251140 1 180 $X=150200 $Y=250780
X41 402 403 11 10 CLKINVX1 $T=154280 251140 0 180 $X=151940 $Y=245320
X42 404 405 11 10 CLKINVX1 $T=156600 272020 1 0 $X=156000 $Y=266200
X43 406 407 11 10 CLKINVX1 $T=160660 282460 0 0 $X=160060 $Y=282100
X44 408 409 11 10 CLKINVX1 $T=167040 292900 0 180 $X=164700 $Y=287080
X45 410 411 11 10 CLKINVX1 $T=171100 282460 0 0 $X=170500 $Y=282100
X46 412 413 11 10 CLKINVX1 $T=173420 230260 1 180 $X=171080 $Y=229900
X47 414 415 11 10 CLKINVX1 $T=174000 198940 1 180 $X=171660 $Y=198580
X48 416 417 11 10 CLKINVX1 $T=174000 313780 0 180 $X=171660 $Y=307960
X49 418 419 11 10 CLKINVX1 $T=177480 282460 0 0 $X=176880 $Y=282100
X50 420 421 11 10 CLKINVX1 $T=178640 334660 0 0 $X=178040 $Y=334300
X51 422 423 11 10 CLKINVX1 $T=183860 198940 1 180 $X=181520 $Y=198580
X52 112 424 11 10 CLKINVX1 $T=185600 188500 1 180 $X=183260 $Y=188140
X53 425 426 11 10 CLKINVX1 $T=186180 334660 1 180 $X=183840 $Y=334300
X54 427 428 11 10 CLKINVX1 $T=186760 272020 0 0 $X=186160 $Y=271660
X55 429 430 11 10 CLKINVX1 $T=195460 345100 1 180 $X=193120 $Y=344740
X56 431 432 11 10 CLKINVX1 $T=194300 272020 0 0 $X=193700 $Y=271660
X57 433 434 11 10 CLKINVX1 $T=196040 303340 1 180 $X=193700 $Y=302980
X58 435 436 11 10 CLKINVX1 $T=194300 324220 0 0 $X=193700 $Y=323860
X59 437 438 11 10 CLKINVX1 $T=198360 198940 1 0 $X=197760 $Y=193120
X60 439 440 11 10 CLKINVX1 $T=200100 198940 1 180 $X=197760 $Y=198580
X61 441 442 11 10 CLKINVX1 $T=200100 345100 0 180 $X=197760 $Y=339280
X62 443 444 11 10 CLKINVX1 $T=201840 198940 1 180 $X=199500 $Y=198580
X63 445 446 11 10 CLKINVX1 $T=203580 303340 0 180 $X=201240 $Y=297520
X64 447 448 11 10 CLKINVX1 $T=204740 272020 0 180 $X=202400 $Y=266200
X65 449 450 11 10 CLKINVX1 $T=204160 345100 1 0 $X=203560 $Y=339280
X66 451 452 11 10 CLKINVX1 $T=207060 334660 1 180 $X=204720 $Y=334300
X67 127 126 11 10 CLKINVX1 $T=212860 188500 1 180 $X=210520 $Y=188140
X68 453 454 11 10 CLKINVX1 $T=212860 209380 0 180 $X=210520 $Y=203560
X69 455 456 11 10 CLKINVX1 $T=213440 334660 0 0 $X=212840 $Y=334300
X70 457 458 11 10 CLKINVX1 $T=213440 345100 0 0 $X=212840 $Y=344740
X71 459 460 11 10 CLKINVX1 $T=218080 282460 1 0 $X=217480 $Y=276640
X72 461 462 11 10 CLKINVX1 $T=219240 334660 0 0 $X=218640 $Y=334300
X73 463 464 11 10 CLKINVX1 $T=222720 209380 1 180 $X=220380 $Y=209020
X74 465 466 11 10 CLKINVX1 $T=223880 209380 0 180 $X=221540 $Y=203560
X75 467 468 11 10 CLKINVX1 $T=226200 198940 0 0 $X=225600 $Y=198580
X76 469 470 11 10 CLKINVX1 $T=227360 230260 0 0 $X=226760 $Y=229900
X77 471 472 11 10 CLKINVX1 $T=229100 292900 1 180 $X=226760 $Y=292540
X78 473 474 11 10 CLKINVX1 $T=227940 198940 0 0 $X=227340 $Y=198580
X79 475 476 11 10 CLKINVX1 $T=230840 230260 1 180 $X=228500 $Y=229900
X80 477 478 11 10 CLKINVX1 $T=230840 240700 0 180 $X=228500 $Y=234880
X81 479 480 11 10 CLKINVX1 $T=230260 282460 1 0 $X=229660 $Y=276640
X82 481 482 11 10 CLKINVX1 $T=230840 219820 1 0 $X=230240 $Y=214000
X83 483 484 11 10 CLKINVX1 $T=232580 303340 0 0 $X=231980 $Y=302980
X84 485 486 11 10 CLKINVX1 $T=241280 292900 0 180 $X=238940 $Y=287080
X85 487 488 11 10 CLKINVX1 $T=244760 230260 0 0 $X=244160 $Y=229900
X86 489 490 11 10 CLKINVX1 $T=255780 230260 1 180 $X=253440 $Y=229900
X87 164 491 11 10 CLKINVX1 $T=266800 198940 0 0 $X=266200 $Y=198580
X88 492 493 11 10 CLKINVX1 $T=272020 230260 1 180 $X=269680 $Y=229900
X89 494 495 11 10 CLKINVX1 $T=273180 272020 0 0 $X=272580 $Y=271660
X90 496 497 11 10 CLKINVX1 $T=278980 251140 1 0 $X=278380 $Y=245320
X91 498 499 11 10 CLKINVX1 $T=283620 198940 1 0 $X=283020 $Y=193120
X92 500 501 11 10 CLKINVX1 $T=283620 209380 0 0 $X=283020 $Y=209020
X93 502 503 11 10 CLKINVX1 $T=294640 219820 0 0 $X=294040 $Y=219460
X94 181 504 11 10 CLKINVX1 $T=295220 188500 0 0 $X=294620 $Y=188140
X95 505 506 11 10 CLKINVX1 $T=295800 219820 1 0 $X=295200 $Y=214000
X96 178 507 11 10 CLKINVX1 $T=299280 198940 0 0 $X=298680 $Y=198580
X97 508 509 11 10 CLKINVX1 $T=301600 198940 0 180 $X=299260 $Y=193120
X98 510 511 11 10 CLKINVX1 $T=303340 198940 1 180 $X=301000 $Y=198580
X99 512 513 11 10 CLKINVX1 $T=303340 209380 0 0 $X=302740 $Y=209020
X100 185 179 11 10 CLKINVX1 $T=307980 188500 1 180 $X=305640 $Y=188140
X101 514 515 11 10 CLKINVX1 $T=306820 219820 1 0 $X=306220 $Y=214000
X102 183 188 11 10 CLKINVX1 $T=307980 188500 0 0 $X=307380 $Y=188140
X103 516 517 11 10 CLKINVX1 $T=310880 198940 1 0 $X=310280 $Y=193120
X104 518 519 11 10 CLKINVX1 $T=312620 198940 1 180 $X=310280 $Y=198580
X105 520 521 11 10 CLKINVX1 $T=313200 261580 1 180 $X=310860 $Y=261220
X106 522 523 11 10 CLKINVX1 $T=316100 209380 1 180 $X=313760 $Y=209020
X107 524 525 11 10 CLKINVX1 $T=319580 198940 0 180 $X=317240 $Y=193120
X108 526 527 11 10 CLKINVX1 $T=327700 261580 1 0 $X=327100 $Y=255760
X109 528 529 11 10 CLKINVX1 $T=328860 240700 0 0 $X=328260 $Y=240340
X110 530 531 11 10 CLKINVX1 $T=330600 313780 0 180 $X=328260 $Y=307960
X111 192 532 11 10 CLKINVX1 $T=330600 198940 1 0 $X=330000 $Y=193120
X112 533 534 11 10 CLKINVX1 $T=339880 365980 0 180 $X=337540 $Y=360160
X113 535 536 11 10 CLKINVX1 $T=342200 345100 0 0 $X=341600 $Y=344740
X114 537 538 11 10 CLKINVX1 $T=343940 272020 1 0 $X=343340 $Y=266200
X115 539 540 11 10 CLKINVX1 $T=348000 251140 0 0 $X=347400 $Y=250780
X116 541 542 11 10 CLKINVX1 $T=350320 303340 1 0 $X=349720 $Y=297520
X117 543 544 11 10 CLKINVX1 $T=353220 240700 0 180 $X=350880 $Y=234880
X118 545 546 11 10 CLKINVX1 $T=353800 230260 1 180 $X=351460 $Y=229900
X119 547 548 11 10 CLKINVX1 $T=359020 261580 1 180 $X=356680 $Y=261220
X120 549 550 11 10 CLKINVX1 $T=358440 251140 1 0 $X=357840 $Y=245320
X121 551 552 11 10 CLKINVX1 $T=360760 261580 0 180 $X=358420 $Y=255760
X122 553 554 11 10 CLKINVX1 $T=360760 334660 1 180 $X=358420 $Y=334300
X123 555 556 11 10 CLKINVX1 $T=360180 209380 0 0 $X=359580 $Y=209020
X124 557 558 11 10 CLKINVX1 $T=361340 198940 1 0 $X=360740 $Y=193120
X125 559 560 11 10 CLKINVX1 $T=363660 313780 0 180 $X=361320 $Y=307960
X126 561 562 11 10 CLKINVX1 $T=368300 230260 0 0 $X=367700 $Y=229900
X127 563 564 11 10 CLKINVX1 $T=368880 355540 0 0 $X=368280 $Y=355180
X128 565 566 11 10 CLKINVX1 $T=371780 251140 0 180 $X=369440 $Y=245320
X129 567 568 11 10 CLKINVX1 $T=371780 240700 0 0 $X=371180 $Y=240340
X130 569 570 11 10 CLKINVX1 $T=374100 240700 0 0 $X=373500 $Y=240340
X131 571 572 11 10 CLKINVX1 $T=380480 355540 1 0 $X=379880 $Y=349720
X132 573 574 11 10 CLKINVX1 $T=386860 303340 1 180 $X=384520 $Y=302980
X133 575 576 11 10 CLKINVX1 $T=392080 240700 1 180 $X=389740 $Y=240340
X134 577 578 11 10 CLKINVX1 $T=393820 272020 0 0 $X=393220 $Y=271660
X135 579 580 11 10 CLKINVX1 $T=394980 324220 0 0 $X=394380 $Y=323860
X136 581 582 11 10 CLKINVX1 $T=397880 240700 1 180 $X=395540 $Y=240340
X137 583 584 11 10 CLKINVX1 $T=397880 261580 1 180 $X=395540 $Y=261220
X138 585 586 11 10 CLKINVX1 $T=397880 240700 0 0 $X=397280 $Y=240340
X139 587 588 11 10 CLKINVX1 $T=399620 303340 1 180 $X=397280 $Y=302980
X140 589 590 11 10 CLKINVX1 $T=399040 292900 0 0 $X=398440 $Y=292540
X141 591 592 11 10 CLKINVX1 $T=401940 355540 0 180 $X=399600 $Y=349720
X142 593 594 11 10 CLKINVX1 $T=402520 292900 1 180 $X=400180 $Y=292540
X143 595 596 11 10 CLKINVX1 $T=403680 324220 0 180 $X=401340 $Y=318400
X144 597 598 11 10 CLKINVX1 $T=402520 355540 0 0 $X=401920 $Y=355180
X145 599 600 11 10 CLKINVX1 $T=406000 355540 1 180 $X=403660 $Y=355180
X146 601 602 11 10 CLKINVX1 $T=408900 261580 0 180 $X=406560 $Y=255760
X147 603 604 11 10 CLKINVX1 $T=408900 292900 1 180 $X=406560 $Y=292540
X148 605 606 11 10 CLKINVX1 $T=408900 313780 0 180 $X=406560 $Y=307960
X149 607 608 11 10 CLKINVX1 $T=410640 324220 0 180 $X=408300 $Y=318400
X150 609 610 11 10 CLKINVX1 $T=410060 303340 0 0 $X=409460 $Y=302980
X151 611 612 11 10 CLKINVX1 $T=410640 198940 0 0 $X=410040 $Y=198580
X152 613 614 11 10 CLKINVX1 $T=413540 324220 0 180 $X=411200 $Y=318400
X153 615 616 11 10 CLKINVX1 $T=414700 272020 0 0 $X=414100 $Y=271660
X154 617 618 11 10 CLKINVX1 $T=416440 365980 0 180 $X=414100 $Y=360160
X155 619 620 11 10 CLKINVX1 $T=419340 355540 1 180 $X=417000 $Y=355180
X156 621 622 11 10 CLKINVX1 $T=419340 313780 1 0 $X=418740 $Y=307960
X157 623 624 11 10 CLKINVX1 $T=424560 345100 0 0 $X=423960 $Y=344740
X158 625 626 11 10 CLKINVX1 $T=429200 355540 0 180 $X=426860 $Y=349720
X159 627 628 11 10 CLKINVX1 $T=429200 365980 1 0 $X=428600 $Y=360160
X160 629 630 11 10 CLKINVX1 $T=432100 219820 0 180 $X=429760 $Y=214000
X161 631 632 11 10 CLKINVX1 $T=431520 261580 1 0 $X=430920 $Y=255760
X162 633 634 11 10 CLKINVX1 $T=432100 282460 0 0 $X=431500 $Y=282100
X163 635 636 11 10 CLKINVX1 $T=433840 292900 0 180 $X=431500 $Y=287080
X164 637 638 11 10 CLKINVX1 $T=436160 345100 1 180 $X=433820 $Y=344740
X165 639 640 11 10 CLKINVX1 $T=437320 292900 1 180 $X=434980 $Y=292540
X166 641 642 11 10 CLKINVX1 $T=437320 365980 0 180 $X=434980 $Y=360160
X167 643 644 11 10 CLKINVX1 $T=436740 251140 0 0 $X=436140 $Y=250780
X168 645 646 11 10 CLKINVX1 $T=437320 292900 0 0 $X=436720 $Y=292540
X169 647 648 11 10 CLKINVX1 $T=438480 251140 0 0 $X=437880 $Y=250780
X170 251 249 11 10 CLKINVX1 $T=442540 376420 0 180 $X=440200 $Y=370600
X171 649 650 11 10 CLKINVX1 $T=441960 324220 1 0 $X=441360 $Y=318400
X172 651 652 11 10 CLKINVX1 $T=445440 251140 0 180 $X=443100 $Y=245320
X173 653 654 11 10 CLKINVX1 $T=446600 303340 1 180 $X=444260 $Y=302980
X174 655 656 11 10 CLKINVX1 $T=446020 355540 0 0 $X=445420 $Y=355180
X175 657 658 11 10 CLKINVX1 $T=446600 282460 1 0 $X=446000 $Y=276640
X176 659 660 11 10 CLKINVX1 $T=447760 313780 0 0 $X=447160 $Y=313420
X177 661 662 11 10 CLKINVX1 $T=447760 334660 1 0 $X=447160 $Y=328840
X178 663 664 11 10 CLKINVX1 $T=448340 261580 1 0 $X=447740 $Y=255760
X179 254 665 11 10 CLKINVX1 $T=450080 198940 0 0 $X=449480 $Y=198580
X180 666 667 11 10 CLKINVX1 $T=452400 209380 1 0 $X=451800 $Y=203560
X181 668 669 11 10 CLKINVX1 $T=455300 355540 1 180 $X=452960 $Y=355180
X182 670 671 11 10 CLKINVX1 $T=454140 376420 1 0 $X=453540 $Y=370600
X183 672 673 11 10 CLKINVX1 $T=454720 313780 0 0 $X=454120 $Y=313420
X184 674 255 11 10 CLKINVX1 $T=457040 188500 1 180 $X=454700 $Y=188140
X185 675 676 11 10 CLKINVX1 $T=458200 345100 1 180 $X=455860 $Y=344740
X186 677 678 11 10 CLKINVX1 $T=457040 376420 1 0 $X=456440 $Y=370600
X187 679 680 11 10 CLKINVX1 $T=457620 240700 1 0 $X=457020 $Y=234880
X188 681 257 11 10 CLKINVX1 $T=459940 188500 1 180 $X=457600 $Y=188140
X189 682 683 11 10 CLKINVX1 $T=458780 240700 0 0 $X=458180 $Y=240340
X190 684 685 11 10 CLKINVX1 $T=458780 251140 0 0 $X=458180 $Y=250780
X191 686 687 11 10 CLKINVX1 $T=460520 324220 0 180 $X=458180 $Y=318400
X192 688 689 11 10 CLKINVX1 $T=459940 272020 0 0 $X=459340 $Y=271660
X193 690 691 11 10 CLKINVX1 $T=460520 292900 1 0 $X=459920 $Y=287080
X194 692 693 11 10 CLKINVX1 $T=460520 324220 1 0 $X=459920 $Y=318400
X195 694 695 11 10 CLKINVX1 $T=464000 324220 1 180 $X=461660 $Y=323860
X196 696 697 11 10 CLKINVX1 $T=462840 313780 0 0 $X=462240 $Y=313420
X197 698 699 11 10 CLKINVX1 $T=465740 355540 0 180 $X=463400 $Y=349720
X198 700 701 11 10 CLKINVX1 $T=469800 313780 1 180 $X=467460 $Y=313420
X199 702 703 11 10 CLKINVX1 $T=468060 355540 0 0 $X=467460 $Y=355180
X200 704 705 11 10 CLKINVX1 $T=471540 313780 1 180 $X=469200 $Y=313420
X201 706 707 11 10 CLKINVX1 $T=470960 272020 1 0 $X=470360 $Y=266200
X202 708 709 11 10 CLKINVX1 $T=471540 251140 0 0 $X=470940 $Y=250780
X203 270 710 11 10 CLKINVX1 $T=473860 198940 0 180 $X=471520 $Y=193120
X204 711 712 11 10 CLKINVX1 $T=475020 240700 0 180 $X=472680 $Y=234880
X205 713 714 11 10 CLKINVX1 $T=475020 240700 1 180 $X=472680 $Y=240340
X206 269 715 11 10 CLKINVX1 $T=476760 198940 0 180 $X=474420 $Y=193120
X207 716 717 11 10 CLKINVX1 $T=478500 240700 1 0 $X=477900 $Y=234880
X208 718 719 11 10 CLKINVX1 $T=483140 240700 0 180 $X=480800 $Y=234880
X209 720 721 11 10 CLKINVX1 $T=481980 251140 1 0 $X=481380 $Y=245320
X210 722 723 11 10 CLKINVX1 $T=483720 324220 1 180 $X=481380 $Y=323860
X211 724 725 11 10 CLKINVX1 $T=484880 334660 0 180 $X=482540 $Y=328840
X212 726 727 11 10 CLKINVX1 $T=485460 355540 1 0 $X=484860 $Y=349720
X213 728 729 11 10 CLKINVX1 $T=487200 324220 0 0 $X=486600 $Y=323860
X214 730 731 11 10 CLKINVX1 $T=487780 251140 0 0 $X=487180 $Y=250780
X215 732 733 11 10 CLKINVX1 $T=491260 251140 1 180 $X=488920 $Y=250780
X216 734 735 11 10 CLKINVX1 $T=490680 324220 1 0 $X=490080 $Y=318400
X217 736 737 11 10 CLKINVX1 $T=496480 230260 1 180 $X=494140 $Y=229900
X218 738 739 11 10 CLKINVX1 $T=504600 230260 1 180 $X=502260 $Y=229900
X219 740 741 11 10 CLKINVX1 $T=504020 251140 1 0 $X=503420 $Y=245320
X220 742 743 11 10 CLKINVX1 $T=505760 334660 1 180 $X=503420 $Y=334300
X221 744 745 11 10 CLKINVX1 $T=506920 240700 0 180 $X=504580 $Y=234880
X222 746 747 11 10 CLKINVX1 $T=510400 345100 0 180 $X=508060 $Y=339280
X223 748 749 11 10 CLKINVX1 $T=510400 334660 1 0 $X=509800 $Y=328840
X224 750 751 11 10 CLKINVX1 $T=513880 324220 0 0 $X=513280 $Y=323860
X225 752 753 11 10 CLKINVX1 $T=519680 240700 0 0 $X=519080 $Y=240340
X226 754 755 11 10 CLKINVX1 $T=520260 261580 1 0 $X=519660 $Y=255760
X227 316 756 11 10 CLKINVX1 $T=531280 198940 0 180 $X=528940 $Y=193120
X228 28 29 11 10 23 330 DFFRHQX1 $T=51040 376420 0 180 $X=34780 $Y=370600
X229 34 29 11 10 23 331 DFFRHQX1 $T=52780 365980 1 180 $X=36520 $Y=365620
X230 757 29 11 10 36 758 DFFRHQX1 $T=54520 303340 1 0 $X=53920 $Y=297520
X231 759 29 11 10 102 760 DFFRHQX1 $T=270280 303340 1 0 $X=269680 $Y=297520
X232 761 29 11 10 221 762 DFFRHQX1 $T=495320 272020 0 180 $X=479060 $Y=266200
X233 268 29 11 10 221 763 DFFRHQX1 $T=485460 365980 1 0 $X=484860 $Y=360160
X234 31 29 11 10 23 42 764 35 SDFFRHQX1 $T=51040 376420 1 0 $X=50440 $Y=370600
X235 765 29 11 10 102 137 766 61 SDFFRHQX1 $T=232580 365980 0 180 $X=212840 $Y=360160
X236 767 11 10 24 29 23 332 DFFRX1 $T=49300 355540 0 0 $X=48700 $Y=355180
X237 768 11 10 769 29 36 770 DFFRX1 $T=52200 282460 0 0 $X=51600 $Y=282100
X238 771 11 10 772 29 36 773 DFFRX1 $T=52780 282460 1 0 $X=52180 $Y=276640
X239 32 11 10 774 29 36 775 DFFRX1 $T=53360 198940 0 0 $X=52760 $Y=198580
X240 26 11 10 776 29 36 777 DFFRX1 $T=53940 209380 1 0 $X=53340 $Y=203560
X241 778 11 10 779 29 36 780 DFFRX1 $T=54520 292900 1 0 $X=53920 $Y=287080
X242 41 11 10 38 29 36 781 DFFRX1 $T=64960 209380 0 0 $X=64360 $Y=209020
X243 782 11 10 783 29 36 784 DFFRX1 $T=64960 230260 0 0 $X=64360 $Y=229900
X244 785 11 10 56 29 36 786 DFFRX1 $T=99760 188500 1 180 $X=82340 $Y=188140
X245 787 11 10 788 29 36 789 DFFRX1 $T=84100 251140 0 0 $X=83500 $Y=250780
X246 790 11 10 791 29 36 792 DFFRX1 $T=84680 272020 1 0 $X=84080 $Y=266200
X247 793 11 10 794 29 36 795 DFFRX1 $T=85260 282460 1 0 $X=84660 $Y=276640
X248 796 11 10 797 29 36 798 DFFRX1 $T=108460 240700 1 0 $X=107860 $Y=234880
X249 799 11 10 800 29 36 801 DFFRX1 $T=108460 240700 0 0 $X=107860 $Y=240340
X250 802 11 10 803 29 36 804 DFFRX1 $T=110780 272020 0 0 $X=110180 $Y=271660
X251 805 11 10 806 29 36 807 DFFRX1 $T=117160 272020 1 0 $X=116560 $Y=266200
X252 808 11 10 809 29 36 810 DFFRX1 $T=125280 240700 0 0 $X=124680 $Y=240340
X253 811 11 10 812 29 36 813 DFFRX1 $T=125860 303340 0 0 $X=125260 $Y=302980
X254 814 11 10 815 29 36 816 DFFRX1 $T=135720 251140 1 0 $X=135120 $Y=245320
X255 817 11 10 818 29 36 819 DFFRX1 $T=153700 230260 0 0 $X=153100 $Y=229900
X256 820 11 10 821 29 36 822 DFFRX1 $T=160080 240700 1 0 $X=159480 $Y=234880
X257 823 11 10 824 29 36 825 DFFRX1 $T=172260 251140 0 0 $X=171660 $Y=250780
X258 826 11 10 827 29 36 828 DFFRX1 $T=175740 251140 1 0 $X=175140 $Y=245320
X259 829 11 10 830 29 36 831 DFFRX1 $T=198360 251140 1 0 $X=197760 $Y=245320
X260 832 11 10 833 29 36 834 DFFRX1 $T=198360 251140 0 0 $X=197760 $Y=250780
X261 835 11 10 836 29 36 837 DFFRX1 $T=215180 251140 1 0 $X=214580 $Y=245320
X262 838 11 10 839 29 36 840 DFFRX1 $T=215180 251140 0 0 $X=214580 $Y=250780
X263 841 11 10 842 29 145 843 DFFRX1 $T=241280 198940 0 180 $X=223860 $Y=193120
X264 844 11 10 845 29 102 846 DFFRX1 $T=227360 240700 0 0 $X=226760 $Y=240340
X265 847 11 10 848 29 102 849 DFFRX1 $T=232000 251140 1 0 $X=231400 $Y=245320
X266 850 11 10 851 29 36 852 DFFRX1 $T=248820 251140 1 180 $X=231400 $Y=250780
X267 853 11 10 162 29 145 155 DFFRX1 $T=256940 188500 1 180 $X=239520 $Y=188140
X268 854 11 10 855 29 145 66 DFFRX1 $T=258100 198940 0 180 $X=240680 $Y=193120
X269 856 11 10 857 29 36 858 DFFRX1 $T=250560 240700 0 0 $X=249960 $Y=240340
X270 859 11 10 860 29 102 861 DFFRX1 $T=270280 209380 1 180 $X=252860 $Y=209020
X271 862 11 10 863 29 36 864 DFFRX1 $T=274920 198940 0 180 $X=257500 $Y=193120
X272 865 11 10 866 29 102 867 DFFRX1 $T=267380 272020 1 0 $X=266780 $Y=266200
X273 868 11 10 869 29 102 870 DFFRX1 $T=269120 261580 1 0 $X=268520 $Y=255760
X274 871 11 10 872 29 102 873 DFFRX1 $T=269120 282460 1 0 $X=268520 $Y=276640
X275 874 11 10 875 29 102 180 DFFRX1 $T=306820 240700 0 180 $X=289400 $Y=234880
X276 876 11 10 877 29 102 878 DFFRX1 $T=307400 240700 1 180 $X=289980 $Y=240340
X277 879 11 10 880 29 102 881 DFFRX1 $T=307980 251140 1 180 $X=290560 $Y=250780
X278 882 11 10 883 29 102 884 DFFRX1 $T=307980 261580 1 180 $X=290560 $Y=261220
X279 885 11 10 886 29 102 887 DFFRX1 $T=305660 251140 1 0 $X=305060 $Y=245320
X280 888 11 10 889 29 102 890 DFFRX1 $T=323640 240700 0 180 $X=306220 $Y=234880
X281 891 11 10 892 29 102 893 DFFRX1 $T=325380 292900 0 180 $X=307960 $Y=287080
X282 894 11 10 895 29 102 896 DFFRX1 $T=309140 240700 0 0 $X=308540 $Y=240340
X283 897 11 10 898 29 193 899 DFFRX1 $T=326540 188500 1 180 $X=309120 $Y=188140
X284 900 11 10 901 29 102 902 DFFRX1 $T=316680 292900 0 0 $X=316080 $Y=292540
X285 903 11 10 904 29 102 905 DFFRX1 $T=341040 251140 0 180 $X=323620 $Y=245320
X286 906 11 10 907 29 102 908 DFFRX1 $T=325380 292900 1 0 $X=324780 $Y=287080
X287 909 11 10 910 29 102 911 DFFRX1 $T=325380 345100 0 0 $X=324780 $Y=344740
X288 201 11 10 912 29 193 196 DFFRX1 $T=343360 188500 1 180 $X=325940 $Y=188140
X289 913 11 10 914 29 102 915 DFFRX1 $T=330600 324220 0 0 $X=330000 $Y=323860
X290 916 11 10 917 29 102 918 DFFRX1 $T=356120 292900 1 180 $X=338700 $Y=292540
X291 919 11 10 920 29 102 921 DFFRX1 $T=342200 292900 1 0 $X=341600 $Y=287080
X292 922 11 10 923 29 193 212 DFFRX1 $T=348000 188500 0 0 $X=347400 $Y=188140
X293 924 11 10 925 29 102 926 DFFRX1 $T=353800 355540 1 0 $X=353200 $Y=349720
X294 927 11 10 928 29 102 929 DFFRX1 $T=354380 324220 0 0 $X=353780 $Y=323860
X295 930 11 10 931 29 102 932 DFFRX1 $T=354380 365980 0 0 $X=353780 $Y=365620
X296 933 11 10 934 29 102 935 DFFRX1 $T=358440 272020 1 0 $X=357840 $Y=266200
X297 936 11 10 937 29 102 938 DFFRX1 $T=359020 292900 1 0 $X=358420 $Y=287080
X298 939 11 10 940 29 102 941 DFFRX1 $T=359020 292900 0 0 $X=358420 $Y=292540
X299 942 11 10 943 29 102 944 DFFRX1 $T=359020 303340 1 0 $X=358420 $Y=297520
X300 945 11 10 946 29 102 947 DFFRX1 $T=378160 324220 0 0 $X=377560 $Y=323860
X301 948 11 10 949 29 221 950 DFFRX1 $T=379320 261580 0 0 $X=378720 $Y=261220
X302 951 11 10 952 29 221 953 DFFRX1 $T=396140 345100 0 180 $X=378720 $Y=339280
X303 954 11 10 955 29 224 956 DFFRX1 $T=396720 230260 0 180 $X=379300 $Y=224440
X304 957 11 10 958 29 224 211 DFFRX1 $T=397300 188500 1 180 $X=379880 $Y=188140
X305 959 11 10 960 29 221 961 DFFRX1 $T=382220 334660 0 0 $X=381620 $Y=334300
X306 962 11 10 963 29 224 964 DFFRX1 $T=402520 230260 1 180 $X=385100 $Y=229900
X307 965 11 10 966 29 221 967 DFFRX1 $T=402520 251140 0 180 $X=385100 $Y=245320
X308 968 11 10 969 29 221 970 DFFRX1 $T=403680 261580 0 180 $X=386260 $Y=255760
X309 971 11 10 972 29 224 202 DFFRX1 $T=412380 209380 1 180 $X=394960 $Y=209020
X310 973 11 10 974 29 221 975 DFFRX1 $T=406000 251140 0 0 $X=405400 $Y=250780
X311 976 11 10 977 29 221 978 DFFRX1 $T=406580 365980 0 0 $X=405980 $Y=365620
X312 979 11 10 980 29 221 981 DFFRX1 $T=433260 272020 1 180 $X=415840 $Y=271660
X313 982 11 10 983 29 221 984 DFFRX1 $T=435580 282460 0 180 $X=418160 $Y=276640
X314 985 11 10 986 29 221 987 DFFRX1 $T=419920 324220 1 0 $X=419320 $Y=318400
X315 988 11 10 989 29 221 990 DFFRX1 $T=420500 313780 0 0 $X=419900 $Y=313420
X316 991 11 10 992 29 224 228 DFFRX1 $T=426300 188500 0 0 $X=425700 $Y=188140
X317 993 11 10 994 29 224 995 DFFRX1 $T=427460 230260 0 0 $X=426860 $Y=229900
X318 996 11 10 997 29 221 998 DFFRX1 $T=429200 240700 0 0 $X=428600 $Y=240340
X319 999 11 10 1000 29 221 1001 DFFRX1 $T=450080 272020 1 180 $X=432660 $Y=271660
X320 1002 11 10 1003 29 221 1004 DFFRX1 $T=459360 334660 1 180 $X=441940 $Y=334300
X321 1005 11 10 1006 29 221 1007 DFFRX1 $T=444280 345100 1 0 $X=443680 $Y=339280
X322 1008 11 10 1009 29 224 1010 DFFRX1 $T=446600 230260 0 0 $X=446000 $Y=229900
X323 1011 11 10 1012 29 221 1013 DFFRX1 $T=446600 303340 0 0 $X=446000 $Y=302980
X324 1014 11 10 261 29 224 253 DFFRX1 $T=465740 219820 1 180 $X=448320 $Y=219460
X325 1015 11 10 1016 29 221 1017 DFFRX1 $T=448920 303340 1 0 $X=448320 $Y=297520
X326 1018 11 10 1019 29 224 277 DFFRX1 $T=468060 209380 0 0 $X=467460 $Y=209020
X327 1020 11 10 1021 29 224 1022 DFFRX1 $T=468060 219820 1 0 $X=467460 $Y=214000
X328 1023 11 10 1024 29 221 1025 DFFRX1 $T=468060 272020 0 0 $X=467460 $Y=271660
X329 1026 11 10 1027 29 221 1028 DFFRX1 $T=484880 345100 0 180 $X=467460 $Y=339280
X330 1029 11 10 1030 29 221 1031 DFFRX1 $T=484880 345100 1 180 $X=467460 $Y=344740
X331 271 11 10 272 29 221 1032 DFFRX1 $T=472120 365980 0 0 $X=471520 $Y=365620
X332 1033 11 10 274 29 224 1034 DFFRX1 $T=499960 188500 1 180 $X=482540 $Y=188140
X333 1035 11 10 1036 29 221 1037 DFFRX1 $T=489520 272020 0 0 $X=488920 $Y=271660
X334 1038 11 10 1039 29 224 285 DFFRX1 $T=507500 209380 0 180 $X=490080 $Y=203560
X335 1040 11 10 1041 29 221 1042 DFFRX1 $T=508080 251140 1 180 $X=490660 $Y=250780
X336 1043 11 10 1044 29 224 244 DFFRX1 $T=510400 219820 0 180 $X=492980 $Y=214000
X337 286 11 10 288 29 221 1045 DFFRX1 $T=493580 365980 0 0 $X=492980 $Y=365620
X338 1046 11 10 1047 29 221 1048 DFFRX1 $T=494740 313780 1 0 $X=494140 $Y=307960
X339 1049 11 10 1050 29 224 1051 DFFRX1 $T=513880 230260 0 180 $X=496460 $Y=224440
X340 1052 11 10 1053 29 221 1054 DFFRX1 $T=498800 272020 1 0 $X=498200 $Y=266200
X341 1055 11 10 1056 29 221 1057 DFFRX1 $T=500540 313780 0 0 $X=499940 $Y=313420
X342 297 11 10 298 29 221 1058 DFFRX1 $T=506340 376420 1 0 $X=505740 $Y=370600
X343 1059 11 10 1060 29 221 1061 DFFRX1 $T=513880 303340 0 0 $X=513280 $Y=302980
X344 1062 11 10 1063 29 221 1064 DFFRX1 $T=515040 313780 1 0 $X=514440 $Y=307960
X345 1065 11 10 1066 29 221 1067 DFFRX1 $T=517360 272020 1 0 $X=516760 $Y=266200
X346 305 11 10 310 29 221 1068 DFFRX1 $T=518520 365980 0 0 $X=517920 $Y=365620
X347 307 11 10 308 29 221 1069 DFFRX1 $T=519100 365980 1 0 $X=518500 $Y=360160
X348 1070 11 10 309 29 221 1071 DFFRX1 $T=519680 355540 0 0 $X=519080 $Y=355180
X349 1072 11 10 1073 29 23 1074 61 58 SDFFRXL $T=80040 365980 0 0 $X=79440 $Y=365620
X350 1075 11 10 1076 29 23 57 61 60 SDFFRXL $T=80620 376420 1 0 $X=80020 $Y=370600
X351 1077 11 10 1078 29 23 1079 61 1080 SDFFRXL $T=108460 334660 0 0 $X=107860 $Y=334300
X352 1081 11 10 1082 29 23 1083 61 1084 SDFFRXL $T=108460 345100 0 0 $X=107860 $Y=344740
X353 1085 11 10 1086 29 23 1087 61 82 SDFFRXL $T=108460 365980 1 0 $X=107860 $Y=360160
X354 1088 11 10 1089 29 23 1090 61 1091 SDFFRXL $T=108460 365980 0 0 $X=107860 $Y=365620
X355 1092 11 10 1093 29 23 1094 61 1095 SDFFRXL $T=109040 345100 1 0 $X=108440 $Y=339280
X356 1096 11 10 1097 29 23 1098 61 1099 SDFFRXL $T=111360 324220 0 0 $X=110760 $Y=323860
X357 1100 11 10 1101 29 23 1102 61 1103 SDFFRXL $T=133400 313780 0 0 $X=132800 $Y=313420
X358 1104 11 10 1105 29 23 1106 61 1107 SDFFRXL $T=135720 324220 0 0 $X=135120 $Y=323860
X359 1108 11 10 1109 29 36 402 1110 403 SDFFRXL $T=142100 240700 0 0 $X=141500 $Y=240340
X360 1111 11 10 1112 29 36 1113 61 1114 SDFFRXL $T=142680 303340 0 0 $X=142080 $Y=302980
X361 1115 11 10 1116 29 23 104 72 105 SDFFRXL $T=147320 376420 1 0 $X=146720 $Y=370600
X362 1117 11 10 1118 29 36 1119 61 1120 SDFFRXL $T=154280 313780 0 0 $X=153680 $Y=313420
X363 1121 11 10 1122 29 102 106 72 103 SDFFRXL $T=154280 365980 0 0 $X=153680 $Y=365620
X364 1123 11 10 1124 29 36 400 1110 401 SDFFRXL $T=175740 251140 0 180 $X=154260 $Y=245320
X365 67 11 10 75 29 36 414 108 415 SDFFRXL $T=157760 198940 1 0 $X=157160 $Y=193120
X366 1125 11 10 1126 29 23 1127 61 1128 SDFFRXL $T=159500 355540 1 0 $X=158900 $Y=349720
X367 1129 11 10 1130 29 23 1131 72 110 SDFFRXL $T=160080 365980 1 0 $X=159480 $Y=360160
X368 1132 11 10 1133 29 36 1134 61 1135 SDFFRXL $T=175160 313780 0 0 $X=174560 $Y=313420
X369 1136 11 10 1137 29 23 1138 61 1139 SDFFRXL $T=175160 324220 1 0 $X=174560 $Y=318400
X370 1140 11 10 1141 29 102 113 72 115 SDFFRXL $T=175160 365980 0 0 $X=174560 $Y=365620
X371 1142 11 10 1143 29 23 1144 61 1145 SDFFRXL $T=198360 313780 1 0 $X=197760 $Y=307960
X372 1146 11 10 1147 29 102 1148 61 1149 SDFFRXL $T=198360 355540 0 0 $X=197760 $Y=355180
X373 1150 11 10 1151 29 102 130 72 132 SDFFRXL $T=198360 365980 0 0 $X=197760 $Y=365620
X374 1152 11 10 1153 29 102 129 72 136 SDFFRXL $T=198360 376420 1 0 $X=197760 $Y=370600
X375 1154 11 10 1155 29 102 1156 61 1157 SDFFRXL $T=203000 303340 0 0 $X=202400 $Y=302980
X376 1158 11 10 1159 29 102 1160 61 1161 SDFFRXL $T=207640 303340 1 0 $X=207040 $Y=297520
X377 1162 11 10 1163 29 102 1164 61 1165 SDFFRXL $T=215180 345100 1 0 $X=214580 $Y=339280
X378 1166 11 10 1167 29 102 140 72 147 SDFFRXL $T=219240 376420 1 0 $X=218640 $Y=370600
X379 1168 11 10 1169 29 102 1170 61 1171 SDFFRXL $T=220980 345100 0 0 $X=220380 $Y=344740
X380 1172 11 10 1173 29 102 1174 61 1175 SDFFRXL $T=228520 303340 1 0 $X=227920 $Y=297520
X381 1176 11 10 1177 29 102 1178 61 1179 SDFFRXL $T=236060 292900 0 0 $X=235460 $Y=292540
X382 1180 11 10 1181 29 102 1182 61 1183 SDFFRXL $T=236060 303340 0 0 $X=235460 $Y=302980
X383 1184 11 10 1185 29 102 1186 61 1187 SDFFRXL $T=256940 345100 0 180 $X=235460 $Y=339280
X384 1188 11 10 1189 29 102 1190 61 1191 SDFFRXL $T=249400 303340 1 0 $X=248800 $Y=297520
X385 1192 11 10 1193 29 102 169 72 171 SDFFRXL $T=263900 376420 1 0 $X=263300 $Y=370600
X386 1194 11 10 1195 29 102 1196 61 1197 SDFFRXL $T=265060 355540 1 0 $X=264460 $Y=349720
X387 1198 11 10 1199 29 102 170 72 173 SDFFRXL $T=265060 355540 0 0 $X=264460 $Y=355180
X388 1200 11 10 1201 29 102 165 61 1202 SDFFRXL $T=265060 365980 1 0 $X=264460 $Y=360160
X389 1203 11 10 1204 29 102 149 61 1205 SDFFRXL $T=265060 365980 0 0 $X=264460 $Y=365620
X390 1206 11 10 1207 29 221 613 608 614 SDFFRXL $T=392080 334660 1 0 $X=391480 $Y=328840
X391 1208 11 10 1209 29 221 595 580 596 SDFFRXL $T=418760 324220 1 180 $X=397280 $Y=323860
X392 1210 11 10 1211 29 224 629 242 630 SDFFRXL $T=448920 219820 1 180 $X=427440 $Y=219460
X393 1212 11 10 1213 29 224 629 1214 630 SDFFRXL $T=449500 230260 0 180 $X=428020 $Y=224440
X394 1215 11 10 1216 29 221 707 1217 706 SDFFRXL $T=488940 261580 1 180 $X=467460 $Y=261220
X395 1218 11 10 1219 29 221 730 733 731 SDFFRXL $T=477340 261580 1 0 $X=476740 $Y=255760
X396 30 32 11 10 1220 44 XNOR3X1 $T=51620 188500 0 0 $X=51020 $Y=188140
X397 783 778 11 10 1221 777 XNOR3X1 $T=52780 219820 1 0 $X=52180 $Y=214000
X398 757 768 11 10 1222 775 XNOR3X1 $T=52780 251140 0 0 $X=52180 $Y=250780
X399 1093 25 11 10 1223 758 XNOR3X1 $T=52780 334660 0 0 $X=52180 $Y=334300
X400 1078 1072 11 10 1224 773 XNOR3X1 $T=59160 334660 1 0 $X=58560 $Y=328840
X401 1093 1100 11 10 1225 784 XNOR3X1 $T=59740 324220 1 0 $X=59140 $Y=318400
X402 794 771 11 10 1226 47 XNOR3X1 $T=63800 251140 1 0 $X=63200 $Y=245320
X403 768 1109 11 10 1227 781 XNOR3X1 $T=66120 219820 0 0 $X=65520 $Y=219460
X404 1078 1112 11 10 1228 770 XNOR3X1 $T=86420 282460 1 180 $X=68420 $Y=282100
X405 782 1109 11 10 1229 50 XNOR3X1 $T=71340 219820 1 0 $X=70740 $Y=214000
X406 793 1109 11 10 1230 52 XNOR3X1 $T=72500 209380 1 0 $X=71900 $Y=203560
X407 776 41 11 10 1231 861 XNOR3X1 $T=73660 198940 0 0 $X=73060 $Y=198580
X408 1082 1075 11 10 1232 780 XNOR3X1 $T=92220 345100 1 180 $X=74220 $Y=344740
X409 788 790 11 10 1233 59 XNOR3X1 $T=86420 251140 1 0 $X=85820 $Y=245320
X410 1097 1112 11 10 1234 795 XNOR3X1 $T=86420 282460 0 0 $X=85820 $Y=282100
X411 1097 1088 11 10 1235 792 XNOR3X1 $T=86420 324220 0 0 $X=85820 $Y=323860
X412 1082 1104 11 10 1236 798 XNOR3X1 $T=108460 303340 0 0 $X=107860 $Y=302980
X413 803 805 11 10 1237 80 XNOR3X1 $T=111940 251140 1 0 $X=111340 $Y=245320
X414 812 1146 11 10 1238 804 XNOR3X1 $T=118900 282460 0 0 $X=118300 $Y=282100
X415 41 75 11 10 86 843 XNOR3X1 $T=119480 198940 1 0 $X=118880 $Y=193120
X416 809 814 11 10 1239 93 XNOR3X1 $T=125280 240700 1 0 $X=124680 $Y=234880
X417 1143 1111 11 10 1240 807 XNOR3X1 $T=145000 272020 1 180 $X=127000 $Y=271660
X418 1130 83 11 10 1241 1103 XNOR3X1 $T=129340 334660 0 0 $X=128740 $Y=334300
X419 1159 1111 11 10 1242 810 XNOR3X1 $T=151380 272020 0 180 $X=133380 $Y=266200
X420 92 67 11 10 95 899 XNOR3X1 $T=137460 188500 0 0 $X=136860 $Y=188140
X421 1130 91 11 10 1243 1102 XNOR3X1 $T=137460 334660 1 0 $X=136860 $Y=328840
X422 30 67 11 10 96 864 XNOR3X1 $T=138620 198940 1 0 $X=138020 $Y=193120
X423 821 796 11 10 1244 101 XNOR3X1 $T=142680 240700 1 0 $X=142080 $Y=234880
X424 818 1109 11 10 1245 97 XNOR3X1 $T=145000 209380 1 0 $X=144400 $Y=203560
X425 1173 1112 11 10 1246 819 XNOR3X1 $T=145000 272020 0 0 $X=144400 $Y=271660
X426 1101 1177 11 10 1247 822 XNOR3X1 $T=152540 251140 0 0 $X=151940 $Y=250780
X427 857 817 11 10 1248 107 XNOR3X1 $T=154280 209380 0 0 $X=153680 $Y=209020
X428 1153 91 11 10 1249 1113 XNOR3X1 $T=172260 313780 0 180 $X=154260 $Y=307960
X429 91 1121 11 10 1250 1120 XNOR3X1 $T=161240 334660 0 0 $X=160640 $Y=334300
X430 1153 1166 11 10 421 1098 XNOR3X1 $T=181540 324220 1 180 $X=163540 $Y=323860
X431 1153 1166 11 10 449 1099 XNOR3X1 $T=181540 334660 0 180 $X=163540 $Y=328840
X432 1126 1117 11 10 1251 825 XNOR3X1 $T=166460 292900 0 0 $X=165860 $Y=292540
X433 1143 1162 11 10 1252 816 XNOR3X1 $T=186760 272020 1 180 $X=168760 $Y=271660
X434 1117 1177 11 10 1253 831 XNOR3X1 $T=173420 261580 0 0 $X=172820 $Y=261220
X435 1137 1132 11 10 1254 834 XNOR3X1 $T=174000 313780 1 0 $X=173400 $Y=307960
X436 1104 1177 11 10 1255 828 XNOR3X1 $T=174580 261580 1 0 $X=173980 $Y=255760
X437 821 1124 11 10 1256 118 XNOR3X1 $T=178640 198940 1 0 $X=178040 $Y=193120
X438 827 823 11 10 1257 117 XNOR3X1 $T=178640 240700 1 0 $X=178040 $Y=234880
X439 833 829 11 10 1258 128 XNOR3X1 $T=198360 209380 0 0 $X=197760 $Y=209020
X440 91 1150 11 10 436 1157 XNOR3X1 $T=198360 324220 0 0 $X=197760 $Y=323860
X441 91 1150 11 10 441 1156 XNOR3X1 $T=198940 324220 1 0 $X=198340 $Y=318400
X442 836 838 11 10 1259 133 XNOR3X1 $T=206480 230260 1 0 $X=205880 $Y=224440
X443 1169 1154 11 10 1260 840 XNOR3X1 $T=206480 292900 1 0 $X=205880 $Y=287080
X444 1193 1153 11 10 1261 1145 XNOR3X1 $T=223880 313780 1 180 $X=205880 $Y=313420
X445 1155 1177 11 10 1262 846 XNOR3X1 $T=218660 261580 0 0 $X=218060 $Y=261220
X446 844 1124 11 10 1263 150 XNOR3X1 $T=222140 188500 0 0 $X=221540 $Y=188140
X447 1199 1153 11 10 1264 1175 XNOR3X1 $T=228520 324220 1 0 $X=227920 $Y=318400
X448 1159 1184 11 10 1265 858 XNOR3X1 $T=233740 272020 0 0 $X=233140 $Y=271660
X449 848 1123 11 10 1266 156 XNOR3X1 $T=236060 209380 0 0 $X=235460 $Y=209020
X450 1173 1180 11 10 1267 849 XNOR3X1 $T=253460 261580 1 180 $X=235460 $Y=261220
X451 868 1124 11 10 1268 158 XNOR3X1 $T=237800 198940 0 0 $X=237200 $Y=198580
X452 848 871 11 10 1269 159 XNOR3X1 $T=239540 230260 1 0 $X=238940 $Y=224440
X453 91 1153 11 10 1270 1179 XNOR3X1 $T=239540 313780 0 0 $X=238940 $Y=313420
X454 91 1152 11 10 1271 1178 XNOR3X1 $T=245920 324220 1 0 $X=245320 $Y=318400
X455 1153 1198 11 10 1272 1174 XNOR3X1 $T=265640 313780 0 180 $X=247640 $Y=307960
X456 1188 1177 11 10 1273 870 XNOR3X1 $T=251140 272020 0 0 $X=250540 $Y=271660
X457 845 865 11 10 1274 166 XNOR3X1 $T=264480 240700 1 0 $X=263880 $Y=234880
X458 759 868 11 10 1275 172 XNOR3X1 $T=267380 240700 0 0 $X=266780 $Y=240340
X459 162 153 11 10 1276 884 XNOR3X1 $T=268540 198940 0 0 $X=267940 $Y=198580
X460 860 862 11 10 1277 878 XNOR3X1 $T=268540 219820 1 0 $X=267940 $Y=214000
X461 1195 1188 11 10 1278 867 XNOR3X1 $T=268540 282460 0 0 $X=267940 $Y=282100
X462 1201 1180 11 10 1279 760 XNOR3X1 $T=268540 313780 1 0 $X=267940 $Y=307960
X463 1204 1184 11 10 1280 873 XNOR3X1 $T=268540 334660 1 0 $X=267940 $Y=328840
X464 862 182 11 10 1281 896 XNOR3X1 $T=301020 219820 0 0 $X=300420 $Y=219460
X465 886 876 11 10 1282 893 XNOR3X1 $T=305080 282460 1 0 $X=304480 $Y=276640
X466 904 882 11 10 1283 902 XNOR3X1 $T=321320 272020 1 0 $X=320720 $Y=266200
X467 889 874 11 10 1284 908 XNOR3X1 $T=323640 240700 1 0 $X=323040 $Y=234880
X468 897 182 11 10 1285 964 XNOR3X1 $T=328280 219820 1 0 $X=327680 $Y=214000
X469 910 1286 11 10 1287 195 XNOR3X1 $T=345680 376420 0 180 $X=327680 $Y=370600
X470 937 906 11 10 1288 911 XNOR3X1 $T=329440 313780 0 0 $X=328840 $Y=313420
X471 914 959 11 10 1289 200 XNOR3X1 $T=329440 334660 1 0 $X=328840 $Y=328840
X472 901 919 11 10 1290 915 XNOR3X1 $T=333500 324220 1 0 $X=332900 $Y=318400
X473 912 182 11 10 203 956 XNOR3X1 $T=334080 198940 1 0 $X=333480 $Y=193120
X474 842 175 11 10 1291 967 XNOR3X1 $T=334080 209380 0 0 $X=333480 $Y=209020
X475 925 1286 11 10 1292 197 XNOR3X1 $T=352060 365980 1 180 $X=334060 $Y=365620
X476 931 1286 11 10 1293 204 XNOR3X1 $T=365980 376420 0 180 $X=347980 $Y=370600
X477 923 210 11 10 1294 935 XNOR3X1 $T=353800 219820 1 0 $X=353200 $Y=214000
X478 943 891 11 10 1295 929 XNOR3X1 $T=371200 324220 0 180 $X=353200 $Y=318400
X479 934 1213 11 10 1296 926 XNOR3X1 $T=356700 282460 0 0 $X=356100 $Y=282100
X480 207 206 11 10 1297 938 XNOR3X1 $T=357280 230260 1 0 $X=356680 $Y=224440
X481 928 1208 11 10 1298 213 XNOR3X1 $T=358440 345100 0 0 $X=357840 $Y=344740
X482 217 219 11 10 1299 950 XNOR3X1 $T=378160 209380 0 0 $X=377560 $Y=209020
X483 895 206 11 10 1300 981 XNOR3X1 $T=378160 251140 0 0 $X=377560 $Y=250780
X484 949 1213 11 10 1301 932 XNOR3X1 $T=395560 282460 0 180 $X=377560 $Y=276640
X485 952 1286 11 10 1302 218 XNOR3X1 $T=395560 376420 0 180 $X=377560 $Y=370600
X486 937 1211 11 10 1303 961 XNOR3X1 $T=381060 324220 1 0 $X=380460 $Y=318400
X487 969 1213 11 10 1304 953 XNOR3X1 $T=399620 282460 1 180 $X=381620 $Y=282100
X488 958 227 11 10 1305 970 XNOR3X1 $T=400780 219820 0 180 $X=382780 $Y=214000
X489 977 1286 11 10 1306 220 XNOR3X1 $T=406580 365980 1 180 $X=388580 $Y=365620
X490 985 1286 11 10 1307 226 XNOR3X1 $T=413540 345100 0 180 $X=395540 $Y=339280
X491 974 1213 11 10 1308 978 XNOR3X1 $T=401360 282460 0 0 $X=400760 $Y=282100
X492 966 208 11 10 1309 984 XNOR3X1 $T=403680 251140 1 0 $X=403080 $Y=245320
X493 232 227 11 10 1310 975 XNOR3X1 $T=405420 209380 1 0 $X=404820 $Y=203560
X494 963 208 11 10 1311 1001 XNOR3X1 $T=406580 230260 0 0 $X=405980 $Y=229900
X495 960 1312 11 10 1313 237 XNOR3X1 $T=407160 345100 0 0 $X=406560 $Y=344740
X496 955 206 11 10 1314 1042 XNOR3X1 $T=409480 219820 0 0 $X=408880 $Y=219460
X497 972 208 11 10 1315 1051 XNOR3X1 $T=412960 219820 1 0 $X=412360 $Y=214000
X498 994 1212 11 10 1316 987 XNOR3X1 $T=419920 261580 0 0 $X=419320 $Y=261220
X499 989 1317 11 10 1318 238 XNOR3X1 $T=439640 345100 0 180 $X=421640 $Y=339280
X500 997 1212 11 10 1319 990 XNOR3X1 $T=422820 251140 1 0 $X=422220 $Y=245320
X501 980 1210 11 10 1320 1004 XNOR3X1 $T=423980 303340 0 0 $X=423380 $Y=302980
X502 240 219 11 10 1321 998 XNOR3X1 $T=428620 209380 1 0 $X=428020 $Y=203560
X503 1011 1286 11 10 1322 234 XNOR3X1 $T=447180 334660 0 180 $X=429180 $Y=328840
X504 992 219 11 10 1323 995 XNOR3X1 $T=433840 219820 1 0 $X=433240 $Y=214000
X505 1009 1212 11 10 1324 1013 XNOR3X1 $T=441380 261580 0 0 $X=440780 $Y=261220
X506 983 1210 11 10 1325 1031 XNOR3X1 $T=443120 292900 1 0 $X=442520 $Y=287080
X507 250 219 11 10 1326 1010 XNOR3X1 $T=444860 209380 0 0 $X=444260 $Y=209020
X508 1000 1210 11 10 1327 1028 XNOR3X1 $T=448340 282460 0 0 $X=447740 $Y=282100
X509 1003 1328 11 10 1329 280 XNOR3X1 $T=468060 365980 1 0 $X=467460 $Y=360160
X510 1024 1218 11 10 1330 763 XNOR3X1 $T=475600 292900 1 0 $X=475000 $Y=287080
X511 1030 1328 11 10 1331 289 XNOR3X1 $T=481400 355540 0 0 $X=480800 $Y=355180
X512 276 1033 11 10 1332 1025 XNOR3X1 $T=500540 198940 1 180 $X=482540 $Y=198580
X513 1036 1286 11 10 1333 1032 XNOR3X1 $T=483720 303340 0 0 $X=483120 $Y=302980
X514 261 1213 11 10 1334 1037 XNOR3X1 $T=486040 240700 0 0 $X=485440 $Y=240340
X515 1026 1312 11 10 1335 295 XNOR3X1 $T=487200 355540 1 0 $X=486600 $Y=349720
X516 1050 1211 11 10 1336 1048 XNOR3X1 $T=493000 261580 0 0 $X=492400 $Y=261220
X517 1036 1052 11 10 1337 1045 XNOR3X1 $T=493580 303340 1 0 $X=492980 $Y=297520
X518 1056 1312 11 10 1338 299 XNOR3X1 $T=498800 355540 0 0 $X=498200 $Y=355180
X519 281 292 11 10 302 1054 XNOR3X1 $T=499960 188500 0 0 $X=499360 $Y=188140
X520 1041 1211 11 10 1339 1057 XNOR3X1 $T=500540 261580 1 0 $X=499940 $Y=255760
X521 1047 1312 11 10 1340 1058 XNOR3X1 $T=505180 355540 1 0 $X=504580 $Y=349720
X522 1044 1211 11 10 1341 1061 XNOR3X1 $T=513880 230260 1 0 $X=513280 $Y=224440
X523 1039 1210 11 10 1342 1064 XNOR3X1 $T=513880 230260 0 0 $X=513280 $Y=229900
X524 1066 1328 11 10 1343 1068 XNOR3X1 $T=516780 303340 1 0 $X=516180 $Y=297520
X525 261 304 11 10 313 1067 XNOR3X1 $T=517360 188500 0 0 $X=516760 $Y=188140
X526 1062 1312 11 10 1344 1069 XNOR3X1 $T=518520 334660 1 0 $X=517920 $Y=328840
X527 1060 1328 11 10 1345 1071 XNOR3X1 $T=519100 345100 1 0 $X=518500 $Y=339280
X528 210 11 10 208 1346 1347 1348 1349 OAI221XL $T=359600 240700 1 0 $X=359000 $Y=234880
X529 1350 11 10 1351 1317 1352 976 571 OAI221XL $T=393240 345100 0 0 $X=392640 $Y=344740
X530 1353 11 10 1354 1212 1355 973 583 OAI221XL $T=411800 261580 0 0 $X=411200 $Y=261220
X531 959 11 10 1328 1356 1357 1358 1359 OAI221XL $T=421660 355540 1 0 $X=421060 $Y=349720
X532 1360 11 10 1361 1317 1362 1035 1363 OAI221XL $T=484300 313780 0 180 $X=477900 $Y=307960
X533 1055 11 10 1328 1364 1365 1366 748 OAI221XL $T=499380 334660 1 0 $X=498780 $Y=328840
X534 1367 11 10 1368 1210 1369 1040 744 OAI221XL $T=512140 240700 1 180 $X=505740 $Y=240340
X535 511 179 11 10 1370 1371 OR3X1 $T=303340 209380 1 180 $X=298100 $Y=209020
X536 540 545 11 10 1372 1373 OR3X1 $T=349740 261580 0 180 $X=344500 $Y=255760
X537 1374 598 11 10 599 1375 OR3X1 $T=406580 355540 0 0 $X=405980 $Y=355180
X538 642 617 11 10 1376 1377 OR3X1 $T=435580 365980 0 180 $X=430340 $Y=360160
X539 723 728 11 10 1378 1379 OR3X1 $T=481980 324220 1 180 $X=476740 $Y=323860
X540 1380 743 11 10 746 1381 OR3X1 $T=504600 345100 0 180 $X=499360 $Y=339280
X541 1382 753 11 10 754 1383 OR3X1 $T=522580 261580 1 180 $X=517340 $Y=261220
X542 793 11 10 1384 1109 351 1385 OAI211XL $T=89900 209380 1 0 $X=89300 $Y=203560
X543 829 11 10 1386 1123 454 1387 OAI211XL $T=202420 209380 0 180 $X=197760 $Y=203560
X544 1388 11 10 1389 421 456 1390 OAI211XL $T=219240 334660 1 180 $X=214580 $Y=334300
X545 844 11 10 138 1124 467 1391 OAI211XL $T=224460 198940 0 180 $X=219800 $Y=193120
X546 862 11 10 1392 182 523 513 OAI211XL $T=309140 209380 1 180 $X=304480 $Y=209020
X547 894 11 10 1393 206 1394 1395 OAI211XL $T=364240 251140 0 180 $X=359580 $Y=245320
X548 979 11 10 1396 1211 635 1397 OAI211XL $T=430360 292900 0 180 $X=425700 $Y=287080
X549 1011 11 10 1398 1286 649 693 OAI211XL $T=444860 313780 1 180 $X=440200 $Y=313420
X550 1008 11 10 1399 1213 679 1400 OAI211XL $T=452400 251140 1 0 $X=451800 $Y=245320
X551 1002 11 10 1401 1312 702 669 OAI211XL $T=459360 355540 1 180 $X=454700 $Y=355180
X552 258 11 10 1402 227 674 262 OAI211XL $T=468060 198940 1 0 $X=467460 $Y=193120
X553 1403 11 10 376 378 77 1404 54 OAI32XL $T=124700 209380 0 0 $X=124100 $Y=209020
X554 98 11 10 405 1405 402 1406 39 OAI32XL $T=156020 261580 1 0 $X=155420 $Y=255760
X555 39 11 10 406 1407 400 1408 98 OAI32XL $T=161240 282460 0 180 $X=155420 $Y=276640
X556 1409 11 10 604 606 595 1410 231 OAI32XL $T=410060 303340 1 180 $X=404240 $Y=302980
X557 1411 11 10 709 721 730 1412 199 OAI32XL $T=482560 251140 0 0 $X=481960 $Y=250780
X558 782 11 10 768 1413 OR2X1 $T=80040 230260 1 0 $X=79440 $Y=224440
X559 1414 11 10 1108 357 OR2X1 $T=88740 219820 1 0 $X=88140 $Y=214000
X560 1108 11 10 783 1415 OR2X1 $T=89320 230260 0 0 $X=88720 $Y=229900
X561 1414 11 10 1109 351 OR2X1 $T=91060 209380 0 0 $X=90460 $Y=209020
X562 788 11 10 794 361 OR2X1 $T=99180 230260 1 0 $X=98580 $Y=224440
X563 55 11 10 785 1416 OR2X1 $T=103240 188500 1 180 $X=99160 $Y=188140
X564 796 11 10 799 1417 OR2X1 $T=104400 240700 0 180 $X=100320 $Y=234880
X565 1418 11 10 1419 65 OR2X1 $T=102660 198940 1 0 $X=102060 $Y=193120
X566 377 11 10 1420 1421 OR2X1 $T=121220 209380 0 0 $X=120620 $Y=209020
X567 1422 11 10 1109 384 OR2X1 $T=129920 209380 0 0 $X=129320 $Y=209020
X568 1423 11 10 1424 1245 OR2X1 $T=135720 209380 1 0 $X=135120 $Y=203560
X569 1109 11 10 818 1425 OR2X1 $T=146160 230260 1 180 $X=142080 $Y=229900
X570 1111 11 10 1143 1426 OR2X1 $T=143840 282460 1 0 $X=143240 $Y=276640
X571 1143 11 10 1159 1427 OR2X1 $T=148480 282460 1 0 $X=147880 $Y=276640
X572 1112 11 10 1173 1428 OR2X1 $T=160080 292900 0 180 $X=156000 $Y=287080
X573 1429 11 10 1177 404 OR2X1 $T=161820 272020 0 180 $X=157740 $Y=266200
X574 91 11 10 1130 1430 OR2X1 $T=161820 324220 1 180 $X=157740 $Y=323860
X575 83 11 10 1121 1431 OR2X1 $T=165300 345100 0 180 $X=161220 $Y=339280
X576 1177 11 10 1101 1432 OR2X1 $T=174000 261580 0 180 $X=169920 $Y=255760
X577 1124 11 10 821 1433 OR2X1 $T=175160 209380 0 0 $X=174560 $Y=209020
X578 1434 11 10 1435 1256 OR2X1 $T=184440 198940 0 0 $X=183840 $Y=198580
X579 1176 11 10 1118 1436 OR2X1 $T=189080 282460 0 0 $X=188480 $Y=282100
X580 1437 11 10 1124 422 OR2X1 $T=194300 209380 0 180 $X=190220 $Y=203560
X581 1438 11 10 1439 1440 OR2X1 $T=196040 198940 1 180 $X=191960 $Y=198580
X582 1150 11 10 91 425 OR2X1 $T=196040 334660 1 180 $X=191960 $Y=334300
X583 83 11 10 1150 429 OR2X1 $T=201840 345100 1 180 $X=197760 $Y=344740
X584 1166 11 10 1153 1390 OR2X1 $T=201840 334660 0 0 $X=201240 $Y=334300
X585 835 11 10 829 1441 OR2X1 $T=202420 209380 1 0 $X=201820 $Y=203560
X586 1152 11 10 1167 1442 OR2X1 $T=205900 345100 1 180 $X=201820 $Y=344740
X587 1152 11 10 1166 457 OR2X1 $T=209960 345100 0 0 $X=209360 $Y=344740
X588 1443 11 10 1444 139 OR2X1 $T=215180 188500 0 0 $X=214580 $Y=188140
X589 836 11 10 845 1445 OR2X1 $T=215180 219820 1 0 $X=214580 $Y=214000
X590 1446 11 10 1123 465 OR2X1 $T=233160 209380 0 180 $X=229080 $Y=203560
X591 1123 11 10 848 1447 OR2X1 $T=232580 209380 0 0 $X=231980 $Y=209020
X592 847 11 10 868 1448 OR2X1 $T=236060 230260 0 180 $X=231980 $Y=224440
X593 1446 11 10 1124 467 OR2X1 $T=237800 198940 1 180 $X=233720 $Y=198580
X594 1153 11 10 1199 1449 OR2X1 $T=242440 324220 0 0 $X=241840 $Y=323860
X595 856 11 10 850 1450 OR2X1 $T=248820 251140 0 0 $X=248220 $Y=250780
X596 841 11 10 854 1451 OR2X1 $T=263320 198940 0 0 $X=262720 $Y=198580
X597 162 11 10 863 516 OR2X1 $T=274920 198940 1 0 $X=274320 $Y=193120
X598 176 11 10 853 1452 OR2X1 $T=289420 188500 0 0 $X=288820 $Y=188140
X599 510 11 10 184 187 OR2X1 $T=302760 188500 0 0 $X=302160 $Y=188140
X600 894 11 10 879 1453 OR2X1 $T=315520 251140 0 0 $X=314920 $Y=250780
X601 842 11 10 898 1454 OR2X1 $T=324220 209380 1 180 $X=320140 $Y=209020
X602 175 11 10 898 1455 OR2X1 $T=326540 209380 0 0 $X=325940 $Y=209020
X603 886 11 10 895 567 OR2X1 $T=338720 240700 0 0 $X=338120 $Y=240340
X604 885 11 10 903 1456 OR2X1 $T=343360 251140 1 0 $X=342760 $Y=245320
X605 539 11 10 1457 1458 OR2X1 $T=348000 240700 0 180 $X=343920 $Y=234880
X606 1459 11 10 206 543 OR2X1 $T=348000 240700 1 0 $X=347400 $Y=234880
X607 1286 11 10 925 1460 OR2X1 $T=349160 345100 0 0 $X=348560 $Y=344740
X608 1213 11 10 934 1461 OR2X1 $T=355540 282460 1 0 $X=354940 $Y=276640
X609 939 11 10 916 1462 OR2X1 $T=359020 303340 0 180 $X=354940 $Y=297520
X610 1459 11 10 208 1349 OR2X1 $T=356120 240700 1 0 $X=355520 $Y=234880
X611 1463 11 10 1464 1297 OR2X1 $T=364820 230260 0 0 $X=364220 $Y=229900
X612 1465 11 10 1317 571 OR2X1 $T=372360 355540 1 0 $X=371760 $Y=349720
X613 1466 11 10 208 569 OR2X1 $T=386860 240700 0 180 $X=382780 $Y=234880
X614 933 11 10 948 1467 OR2X1 $T=383380 272020 1 0 $X=382780 $Y=266200
X615 1465 11 10 1286 597 OR2X1 $T=383380 355540 1 0 $X=382780 $Y=349720
X616 1466 11 10 206 1394 OR2X1 $T=390340 240700 0 180 $X=386260 $Y=234880
X617 1468 11 10 1211 589 OR2X1 $T=388600 292900 0 0 $X=388000 $Y=292540
X618 1468 11 10 1210 1469 OR2X1 $T=389760 303340 1 0 $X=389160 $Y=297520
X619 962 11 10 965 575 OR2X1 $T=396140 240700 1 180 $X=392060 $Y=240340
X620 1470 11 10 1212 583 OR2X1 $T=394400 272020 1 0 $X=393800 $Y=266200
X621 1471 11 10 1472 1303 OR2X1 $T=397880 313780 1 180 $X=393800 $Y=313420
X622 1473 11 10 1474 1306 OR2X1 $T=397880 355540 1 180 $X=393800 $Y=355180
X623 1470 11 10 1213 1475 OR2X1 $T=397300 272020 0 0 $X=396700 $Y=271660
X624 605 11 10 1476 1477 OR2X1 $T=401360 313780 1 180 $X=397280 $Y=313420
X625 208 11 10 963 1478 OR2X1 $T=399040 240700 1 0 $X=398440 $Y=234880
X626 1352 11 10 591 623 OR2X1 $T=400200 345100 0 0 $X=399600 $Y=344740
X627 971 11 10 206 1479 OR2X1 $T=404260 219820 0 180 $X=400180 $Y=214000
X628 968 11 10 1213 1480 OR2X1 $T=406580 272020 0 0 $X=405980 $Y=271660
X629 1481 11 10 1482 1308 OR2X1 $T=412380 282460 1 0 $X=411780 $Y=276640
X630 940 11 10 980 1483 OR2X1 $T=412380 292900 0 0 $X=411780 $Y=292540
X631 1484 11 10 1485 613 OR2X1 $T=412960 313780 0 0 $X=412360 $Y=313420
X632 1486 11 10 1487 1313 OR2X1 $T=412960 355540 1 0 $X=412360 $Y=349720
X633 1488 11 10 611 1489 OR2X1 $T=419340 198940 0 180 $X=415260 $Y=193120
X634 1355 11 10 601 643 OR2X1 $T=416440 261580 1 0 $X=415840 $Y=255760
X635 1209 11 10 1207 1490 OR2X1 $T=418760 345100 1 0 $X=418160 $Y=339280
X636 206 11 10 955 1491 OR2X1 $T=424560 230260 0 180 $X=420480 $Y=224440
X637 1212 11 10 994 1492 OR2X1 $T=421660 261580 1 0 $X=421060 $Y=255760
X638 227 11 10 232 1493 OR2X1 $T=426300 209380 0 180 $X=422220 $Y=203560
X639 1317 11 10 986 1494 OR2X1 $T=430940 324220 1 180 $X=426860 $Y=323860
X640 219 11 10 992 1495 OR2X1 $T=430360 198940 0 0 $X=429760 $Y=198580
X641 1496 11 10 1211 635 OR2X1 $T=436160 282460 0 0 $X=435560 $Y=282100
X642 1496 11 10 1210 639 OR2X1 $T=436160 292900 1 0 $X=435560 $Y=287080
X643 641 11 10 1497 1498 OR2X1 $T=440220 355540 1 180 $X=436140 $Y=355180
X644 1499 11 10 1286 649 OR2X1 $T=437900 324220 1 0 $X=437300 $Y=318400
X645 999 11 10 982 657 OR2X1 $T=439060 282460 1 0 $X=438460 $Y=276640
X646 1206 11 10 1005 1500 OR2X1 $T=440220 345100 1 0 $X=439620 $Y=339280
X647 1016 11 10 1012 672 OR2X1 $T=441380 303340 0 0 $X=440780 $Y=302980
X648 1499 11 10 1317 659 OR2X1 $T=444280 324220 1 0 $X=443680 $Y=318400
X649 1501 11 10 219 254 OR2X1 $T=446600 188500 0 0 $X=446000 $Y=188140
X650 1502 11 10 1212 682 OR2X1 $T=447180 240700 1 0 $X=446580 $Y=234880
X651 1210 11 10 1000 1503 OR2X1 $T=448920 282460 1 0 $X=448320 $Y=276640
X652 1501 11 10 227 674 OR2X1 $T=451240 188500 0 0 $X=450640 $Y=188140
X653 1003 11 10 1006 1504 OR2X1 $T=454720 345100 1 180 $X=450640 $Y=344740
X654 1502 11 10 1213 679 OR2X1 $T=452400 240700 1 0 $X=451800 $Y=234880
X655 1021 11 10 1009 1505 OR2X1 $T=471540 240700 0 180 $X=467460 $Y=234880
X656 1506 11 10 1507 1217 OR2X1 $T=472700 261580 0 180 $X=468620 $Y=255760
X657 1015 11 10 1215 1508 OR2X1 $T=469220 303340 0 0 $X=468620 $Y=302980
X658 1328 11 10 1027 1509 OR2X1 $T=471540 334660 0 0 $X=470940 $Y=334300
X659 1510 11 10 1328 698 OR2X1 $T=477920 355540 1 180 $X=473840 $Y=355180
X660 1511 11 10 1213 711 OR2X1 $T=478500 240700 0 180 $X=474420 $Y=234880
X661 1219 11 10 1216 1512 OR2X1 $T=475020 292900 0 0 $X=474420 $Y=292540
X662 1511 11 10 1212 1513 OR2X1 $T=476760 230260 0 0 $X=476160 $Y=229900
X663 1510 11 10 1312 702 OR2X1 $T=481400 355540 1 180 $X=477320 $Y=355180
X664 720 11 10 1514 1515 OR2X1 $T=483720 251140 1 0 $X=483120 $Y=245320
X665 722 11 10 1516 1517 OR2X1 $T=483720 324220 0 0 $X=483120 $Y=323860
X666 1518 11 10 1519 1333 OR2X1 $T=490680 313780 1 0 $X=490080 $Y=307960
X667 1520 11 10 1521 1334 OR2X1 $T=493000 240700 1 0 $X=492400 $Y=234880
X668 1328 11 10 1046 1522 OR2X1 $T=493580 324220 0 0 $X=492980 $Y=323860
X669 1369 11 10 740 688 OR2X1 $T=504020 251140 0 180 $X=499940 $Y=245320
X670 286 11 10 245 294 OR2X1 $T=502860 376420 1 0 $X=502260 $Y=370600
X671 1523 11 10 1210 744 OR2X1 $T=511560 240700 0 180 $X=507480 $Y=234880
X672 1524 11 10 1525 1338 OR2X1 $T=513880 334660 1 180 $X=509800 $Y=334300
X673 1062 11 10 1059 1526 OR2X1 $T=515040 313780 0 180 $X=510960 $Y=307960
X674 1038 11 10 1043 1527 OR2X1 $T=512140 219820 1 0 $X=511540 $Y=214000
X675 1523 11 10 1211 752 OR2X1 $T=512720 240700 1 0 $X=512120 $Y=234880
X676 1528 11 10 1529 1339 OR2X1 $T=514460 251140 1 0 $X=513860 $Y=245320
X677 1530 11 10 1312 742 OR2X1 $T=519100 334660 1 180 $X=515020 $Y=334300
X678 307 11 10 1070 311 OR2X1 $T=526640 376420 0 180 $X=522560 $Y=370600
X679 1328 11 10 1063 1531 OR2X1 $T=528380 313780 1 180 $X=524300 $Y=313420
X680 1530 11 10 1328 748 OR2X1 $T=529540 334660 1 180 $X=525460 $Y=334300
X681 1414 783 11 10 768 NOR2BXL $T=88160 219820 1 180 $X=84080 $Y=219460
X682 335 800 11 10 797 NOR2BXL $T=97440 230260 0 0 $X=96840 $Y=229900
X683 1532 1125 11 10 1086 NOR2BXL $T=103820 345100 1 180 $X=99740 $Y=344740
X684 1533 1086 11 10 1126 NOR2BXL $T=102080 355540 1 0 $X=101480 $Y=349720
X685 371 787 11 10 806 NOR2BXL $T=108460 219820 1 0 $X=107860 $Y=214000
X686 1422 809 11 10 805 NOR2BXL $T=117160 230260 0 180 $X=113080 $Y=224440
X687 375 37 11 10 1534 NOR2BXL $T=117740 209380 0 0 $X=117140 $Y=209020
X688 373 811 11 10 1097 NOR2BXL $T=118900 292900 0 0 $X=118300 $Y=292540
X689 1535 1112 11 10 1097 NOR2BXL $T=124120 292900 0 180 $X=120040 $Y=287080
X690 1241 1536 11 10 1537 NOR2BXL $T=142680 345100 0 180 $X=138600 $Y=339280
X691 1538 1422 11 10 1109 NOR2BXL $T=145000 209380 0 0 $X=144400 $Y=209020
X692 1539 91 11 10 1130 NOR2BXL $T=150220 334660 0 0 $X=149620 $Y=334300
X693 406 1112 11 10 1427 NOR2BXL $T=154860 282460 1 180 $X=150780 $Y=282100
X694 1540 83 11 10 1130 NOR2BXL $T=160660 334660 1 180 $X=156580 $Y=334300
X695 1541 1542 11 10 1543 NOR2BXL $T=160660 345100 1 180 $X=156580 $Y=344740
X696 1429 1118 11 10 1104 NOR2BXL $T=162400 272020 0 0 $X=161800 $Y=271660
X697 1544 1429 11 10 1177 NOR2BXL $T=165880 272020 0 0 $X=165280 $Y=271660
X698 1545 1122 11 10 83 NOR2BXL $T=165880 345100 0 0 $X=165280 $Y=344740
X699 427 1117 11 10 1105 NOR2BXL $T=167620 282460 0 0 $X=167020 $Y=282100
X700 408 1158 11 10 1143 NOR2BXL $T=183860 292900 0 0 $X=183260 $Y=292540
X701 1546 1437 11 10 1124 NOR2BXL $T=189080 209380 0 0 $X=188480 $Y=209020
X702 1547 1151 11 10 83 NOR2BXL $T=194880 355540 0 180 $X=190800 $Y=349720
X703 1437 827 11 10 829 NOR2BXL $T=192560 209380 0 0 $X=191960 $Y=209020
X704 1548 1151 11 10 91 NOR2BXL $T=198360 334660 0 0 $X=197760 $Y=334300
X705 439 443 11 10 37 NOR2BXL $T=201840 198940 0 0 $X=201240 $Y=198580
X706 1549 1167 11 10 1152 NOR2BXL $T=206480 345100 0 0 $X=205880 $Y=344740
X707 459 1154 11 10 1133 NOR2BXL $T=207640 282460 1 0 $X=207040 $Y=276640
X708 1550 1176 11 10 1155 NOR2BXL $T=211120 282460 1 0 $X=210520 $Y=276640
X709 1551 1193 11 10 1152 NOR2BXL $T=219820 324220 0 180 $X=215740 $Y=318400
X710 1552 765 11 10 1163 NOR2BXL $T=233740 334660 1 180 $X=229660 $Y=334300
X711 1553 1162 11 10 765 NOR2BXL $T=237220 334660 1 180 $X=233140 $Y=334300
X712 1446 848 11 10 868 NOR2BXL $T=234320 209380 1 0 $X=233720 $Y=203560
X713 487 851 11 10 857 NOR2BXL $T=240700 230260 1 180 $X=236620 $Y=229900
X714 1554 1261 11 10 1555 NOR2BXL $T=240700 334660 0 180 $X=236620 $Y=328840
X715 1556 1152 11 10 1199 NOR2BXL $T=248820 334660 1 0 $X=248220 $Y=328840
X716 1557 1558 11 10 1389 NOR2BXL $T=255780 334660 0 180 $X=251700 $Y=328840
X717 500 855 11 10 842 NOR2BXL $T=256940 209380 0 180 $X=252860 $Y=203560
X718 1559 1153 11 10 1199 NOR2BXL $T=261000 334660 1 0 $X=260400 $Y=328840
X719 1272 1557 11 10 1560 NOR2BXL $T=263320 324220 1 0 $X=262720 $Y=318400
X720 1561 183 11 10 1562 NOR2BXL $T=298700 198940 1 180 $X=294620 $Y=198580
X721 520 880 11 10 895 NOR2BXL $T=314360 251140 1 180 $X=310280 $Y=250780
X722 522 182 11 10 1454 NOR2BXL $T=316100 209380 0 0 $X=315500 $Y=209020
X723 1563 897 11 10 842 NOR2BXL $T=324800 198940 1 0 $X=324200 $Y=193120
X724 1459 904 11 10 888 NOR2BXL $T=344520 240700 0 180 $X=340440 $Y=234880
X725 205 182 11 10 201 NOR2BXL $T=346840 188500 1 180 $X=342760 $Y=188140
X726 563 930 11 10 925 NOR2BXL $T=354960 355540 1 180 $X=350880 $Y=355180
X727 1348 206 11 10 210 NOR2BXL $T=359020 230260 1 180 $X=354940 $Y=229900
X728 1465 931 11 10 924 NOR2BXL $T=363660 355540 1 180 $X=359580 $Y=355180
X729 1564 562 11 10 1565 NOR2BXL $T=366560 251140 1 180 $X=362480 $Y=250780
X730 559 917 11 10 940 NOR2BXL $T=364820 313780 1 0 $X=364220 $Y=307960
X731 1566 1206 11 10 946 NOR2BXL $T=375260 334660 1 180 $X=371180 $Y=334300
X732 1567 946 11 10 1207 NOR2BXL $T=378740 334660 0 0 $X=378140 $Y=334300
X733 609 942 11 10 940 NOR2BXL $T=384540 303340 0 180 $X=380460 $Y=297520
X734 1468 943 11 10 919 NOR2BXL $T=389180 303340 0 180 $X=385100 $Y=297520
X735 1470 949 11 10 933 NOR2BXL $T=390340 272020 0 180 $X=386260 $Y=266200
X736 1466 963 11 10 965 NOR2BXL $T=390340 240700 1 0 $X=389740 $Y=234880
X737 585 1568 11 10 1479 NOR2BXL $T=396720 230260 1 0 $X=396120 $Y=224440
X738 591 1317 11 10 952 NOR2BXL $T=405420 355540 0 180 $X=401340 $Y=349720
X739 601 1212 11 10 969 NOR2BXL $T=407160 261580 0 180 $X=403080 $Y=255760
X740 1350 1286 11 10 976 NOR2BXL $T=403680 345100 0 0 $X=403080 $Y=344740
X741 1569 208 11 10 972 NOR2BXL $T=407740 219820 0 180 $X=403660 $Y=214000
X742 599 1286 11 10 952 NOR2BXL $T=406000 355540 1 0 $X=405400 $Y=349720
X743 611 227 11 10 958 NOR2BXL $T=410640 198940 0 180 $X=406560 $Y=193120
X744 1570 219 11 10 958 NOR2BXL $T=410640 198940 1 180 $X=406560 $Y=198580
X745 603 593 11 10 231 NOR2BXL $T=412380 292900 1 180 $X=408300 $Y=292540
X746 1358 1312 11 10 959 NOR2BXL $T=412960 355540 0 180 $X=408880 $Y=349720
X747 1353 1213 11 10 973 NOR2BXL $T=411800 261580 1 0 $X=411200 $Y=255760
X748 1499 986 11 10 988 NOR2BXL $T=418760 324220 0 180 $X=414680 $Y=318400
X749 619 1312 11 10 1490 NOR2BXL $T=419340 355540 0 0 $X=418740 $Y=355180
X750 1502 997 11 10 993 NOR2BXL $T=427460 230260 1 180 $X=423380 $Y=229900
X751 647 996 11 10 994 NOR2BXL $T=428620 251140 1 180 $X=424540 $Y=250780
X752 1571 991 11 10 240 NOR2BXL $T=430360 198940 1 180 $X=426280 $Y=198580
X753 1572 985 11 10 989 NOR2BXL $T=429780 334660 0 0 $X=429180 $Y=334300
X754 1496 1000 11 10 982 NOR2BXL $T=435580 282460 1 0 $X=434980 $Y=276640
X755 1501 992 11 10 247 NOR2BXL $T=446600 188500 1 180 $X=442520 $Y=188140
X756 1573 625 11 10 1574 NOR2BXL $T=445440 355540 1 0 $X=444840 $Y=349720
X757 1575 252 11 10 264 NOR2BXL $T=460520 188500 0 0 $X=459920 $Y=188140
X758 1576 701 11 10 1577 NOR2BXL $T=465740 324220 0 180 $X=461660 $Y=318400
X759 708 716 11 10 199 NOR2BXL $T=471540 251140 1 180 $X=467460 $Y=250780
X760 1578 761 11 10 1216 NOR2BXL $T=474440 292900 0 180 $X=470360 $Y=287080
X761 713 1020 11 10 274 NOR2BXL $T=478500 251140 1 0 $X=477900 $Y=245320
X762 1510 1030 11 10 1026 NOR2BXL $T=481980 355540 0 180 $X=477900 $Y=349720
X763 1579 1215 11 10 761 NOR2BXL $T=484300 292900 1 180 $X=480220 $Y=292540
X764 726 1029 11 10 1027 NOR2BXL $T=485460 355540 0 180 $X=481380 $Y=349720
X765 1511 274 11 10 279 NOR2BXL $T=483140 240700 1 0 $X=482540 $Y=234880
X766 278 1019 11 10 1021 NOR2BXL $T=484880 209380 0 0 $X=484280 $Y=209020
X767 1580 1020 11 10 1019 NOR2BXL $T=484880 219820 1 0 $X=484280 $Y=214000
X768 734 1286 11 10 1512 NOR2BXL $T=488360 303340 0 180 $X=484280 $Y=297520
X769 1360 1286 11 10 1035 NOR2BXL $T=486040 313780 1 0 $X=485440 $Y=307960
X770 1366 1312 11 10 1055 NOR2BXL $T=499380 334660 0 180 $X=495300 $Y=328840
X771 740 1210 11 10 1050 NOR2BXL $T=499960 251140 0 180 $X=495880 $Y=245320
X772 1581 1365 11 10 1522 NOR2BXL $T=501120 324220 1 180 $X=497040 $Y=323860
X773 1523 1044 11 10 1038 NOR2BXL $T=508080 219820 1 180 $X=504000 $Y=219460
X774 746 1312 11 10 1047 NOR2BXL $T=505180 345100 1 0 $X=504580 $Y=339280
X775 1367 1211 11 10 1040 NOR2BXL $T=509240 251140 0 180 $X=505160 $Y=245320
X776 754 1211 11 10 1050 NOR2BXL $T=515620 261580 1 180 $X=511540 $Y=261220
X777 1530 1060 11 10 1062 NOR2BXL $T=520260 334660 0 0 $X=519660 $Y=334300
X778 315 314 11 10 294 NOR2BXL $T=530120 376420 0 180 $X=526040 $Y=370600
X779 1109 362 11 10 351 1534 OA21X1 $T=98600 209380 0 0 $X=98000 $Y=209020
X780 1582 1385 11 10 375 1419 OA21X1 $T=106140 209380 0 180 $X=100320 $Y=203560
X781 388 1583 11 10 37 1418 OA21X1 $T=106140 219820 0 180 $X=100320 $Y=214000
X782 788 1109 11 10 1584 1583 OA21X1 $T=113680 230260 0 180 $X=107860 $Y=224440
X783 1109 371 11 10 1584 1585 OA21X1 $T=111940 219820 1 0 $X=111340 $Y=214000
X784 1111 373 11 10 359 1586 OA21X1 $T=113680 292900 0 0 $X=113080 $Y=292540
X785 809 1109 11 10 1585 1587 OA21X1 $T=130500 219820 1 0 $X=129900 $Y=214000
X786 1116 1122 11 10 83 1536 OA21X1 $T=135140 355540 1 0 $X=134540 $Y=349720
X787 1545 1542 11 10 1431 1588 OA21X1 $T=165880 345100 1 180 $X=160060 $Y=344740
X788 1548 436 11 10 425 1589 OA21X1 $T=194300 324220 1 180 $X=188480 $Y=323860
X789 1547 442 11 10 429 1590 OA21X1 $T=195460 345100 0 180 $X=189640 $Y=339280
X790 1177 459 11 10 1591 1592 OA21X1 $T=198360 261580 0 0 $X=197760 $Y=261220
X791 1593 1391 11 10 439 1444 OA21X1 $T=211120 198940 0 180 $X=205300 $Y=193120
X792 1549 450 11 10 457 1594 OA21X1 $T=205900 345100 1 0 $X=205300 $Y=339280
X793 1166 134 11 10 1153 1388 OA21X1 $T=214020 355540 1 0 $X=213420 $Y=349720
X794 453 1595 11 10 54 1443 OA21X1 $T=215760 198940 0 0 $X=215160 $Y=198580
X795 836 1124 11 10 464 1595 OA21X1 $T=220980 209380 1 180 $X=215160 $Y=209020
X796 1551 1261 11 10 1596 1597 OA21X1 $T=219820 324220 1 0 $X=219220 $Y=318400
X797 1192 163 11 10 1153 1558 OA21X1 $T=257520 334660 1 180 $X=251700 $Y=334300
X798 1199 1152 11 10 1557 1598 OA21X1 $T=255780 334660 1 0 $X=255180 $Y=328840
X799 182 517 11 10 523 185 OA21X1 $T=310880 198940 1 180 $X=305060 $Y=198580
X800 863 175 11 10 1599 512 OA21X1 $T=314360 209380 1 180 $X=308540 $Y=209020
X801 863 182 11 10 524 508 OA21X1 $T=317840 198940 0 180 $X=312020 $Y=193120
X802 182 1563 11 10 192 524 OA21X1 $T=324800 198940 0 180 $X=318980 $Y=193120
X803 175 1563 11 10 194 1599 OA21X1 $T=325960 209380 0 180 $X=320140 $Y=203560
X804 1286 563 11 10 1600 1601 OA21X1 $T=363660 355540 0 0 $X=363060 $Y=355180
X805 568 208 11 10 569 561 OA21X1 $T=375840 240700 0 180 $X=370020 $Y=234880
X806 895 206 11 10 1602 565 OA21X1 $T=378740 251140 1 0 $X=378140 $Y=245320
X807 206 576 11 10 582 1602 OA21X1 $T=390340 240700 1 180 $X=384520 $Y=240340
X808 920 1211 11 10 1603 573 OA21X1 $T=394400 303340 1 0 $X=393800 $Y=297520
X809 958 227 11 10 1604 1605 OA21X1 $T=400200 209380 1 0 $X=399600 $Y=203560
X810 1211 609 11 10 1606 1603 OA21X1 $T=411800 303340 0 180 $X=405980 $Y=297520
X811 940 1211 11 10 1606 1607 OA21X1 $T=411800 303340 1 0 $X=411200 $Y=297520
X812 587 1607 11 10 199 1484 OA21X1 $T=418180 303340 1 180 $X=412360 $Y=302980
X813 1608 1397 11 10 603 1485 OA21X1 $T=419340 313780 0 180 $X=413520 $Y=307960
X814 980 1211 11 10 645 1606 OA21X1 $T=421080 292900 1 0 $X=420480 $Y=287080
X815 1317 1572 11 10 1375 1609 OA21X1 $T=432100 324220 0 0 $X=431500 $Y=323860
X816 1286 1572 11 10 623 661 OA21X1 $T=435000 334660 0 0 $X=434400 $Y=334300
X817 1213 647 11 10 643 651 OA21X1 $T=440220 251140 0 0 $X=439620 $Y=250780
X818 1009 1213 11 10 651 1610 OA21X1 $T=447760 240700 0 0 $X=447160 $Y=240340
X819 219 1571 11 10 1489 1611 OA21X1 $T=448340 198940 1 0 $X=447740 $Y=193120
X820 1012 1286 11 10 661 696 OA21X1 $T=448340 324220 1 0 $X=447740 $Y=318400
X821 1211 658 11 10 688 645 OA21X1 $T=455300 272020 1 180 $X=449480 $Y=271660
X822 1012 1317 11 10 1609 692 OA21X1 $T=450660 324220 0 0 $X=450060 $Y=323860
X823 250 227 11 10 666 681 OA21X1 $T=455300 209380 1 0 $X=454700 $Y=203560
X824 673 1317 11 10 659 700 OA21X1 $T=457040 313780 0 0 $X=456440 $Y=313420
X825 1612 1400 11 10 708 1507 OA21X1 $T=460520 251140 0 0 $X=459920 $Y=250780
X826 1003 1328 11 10 1613 668 OA21X1 $T=465740 355540 1 180 $X=459920 $Y=355180
X827 1021 1213 11 10 1610 1614 OA21X1 $T=473280 240700 1 180 $X=467460 $Y=240340
X828 718 1614 11 10 231 1506 OA21X1 $T=468060 251140 1 0 $X=467460 $Y=245320
X829 1328 726 11 10 1381 1613 OA21X1 $T=478500 355540 0 180 $X=472680 $Y=349720
X830 1213 713 11 10 1610 1615 OA21X1 $T=475020 240700 0 0 $X=474420 $Y=240340
X831 281 1213 11 10 1615 736 OA21X1 $T=488360 219820 1 0 $X=487760 $Y=214000
X832 1417 1221 11 10 37 336 MXI2XL $T=65540 219820 1 180 $X=60300 $Y=219460
X833 334 1222 11 10 37 1616 MXI2XL $T=63220 240700 0 0 $X=62620 $Y=240340
X834 1617 1223 11 10 39 337 MXI2XL $T=68440 345100 1 180 $X=63200 $Y=344740
X835 340 1220 11 10 45 46 MXI2XL $T=73660 188500 1 180 $X=68420 $Y=188140
X836 348 1224 11 10 39 343 MXI2XL $T=74820 334660 1 180 $X=69580 $Y=334300
X837 345 1226 11 10 37 342 MXI2XL $T=71340 251140 0 0 $X=70740 $Y=250780
X838 1618 1228 11 10 39 349 MXI2XL $T=72500 303340 1 0 $X=71900 $Y=297520
X839 1416 1231 11 10 45 51 MXI2XL $T=82940 188500 1 180 $X=77700 $Y=188140
X840 1619 1229 11 10 37 1620 MXI2XL $T=90480 230260 0 180 $X=85240 $Y=224440
X841 1621 1225 11 10 39 1622 MXI2XL $T=90480 313780 0 0 $X=89880 $Y=313420
X842 360 1234 11 10 39 363 MXI2XL $T=91640 292900 0 0 $X=91040 $Y=292540
X843 365 1235 11 10 39 369 MXI2XL $T=96860 334660 0 180 $X=91620 $Y=328840
X844 1623 1233 11 10 37 1624 MXI2XL $T=101500 251140 0 0 $X=100900 $Y=250780
X845 1625 1238 11 10 39 380 MXI2XL $T=131080 292900 1 180 $X=125840 $Y=292540
X846 392 1236 11 10 39 383 MXI2XL $T=127020 313780 0 0 $X=126420 $Y=313420
X847 1626 1239 11 10 37 390 MXI2XL $T=135720 251140 0 180 $X=130480 $Y=245320
X848 387 1240 11 10 39 1627 MXI2XL $T=136300 282460 0 0 $X=135700 $Y=282100
X849 394 1244 11 10 37 399 MXI2XL $T=152540 230260 1 180 $X=147300 $Y=229900
X850 397 1248 11 10 37 1628 MXI2XL $T=148480 209380 0 0 $X=147880 $Y=209020
X851 411 1252 11 10 39 418 MXI2XL $T=172840 282460 0 0 $X=172240 $Y=282100
X852 416 1251 11 10 39 1629 MXI2XL $T=183280 303340 0 180 $X=178040 $Y=297520
X853 412 1257 11 10 37 1630 MXI2XL $T=189660 230260 0 0 $X=189060 $Y=229900
X854 1631 1253 11 10 39 432 MXI2XL $T=198360 272020 1 0 $X=197760 $Y=266200
X855 433 1254 11 10 39 445 MXI2XL $T=198360 303340 0 0 $X=197760 $Y=302980
X856 483 1260 11 10 39 471 MXI2XL $T=228520 292900 0 180 $X=223280 $Y=287080
X857 477 1258 11 10 37 470 MXI2XL $T=225620 230260 1 0 $X=225020 $Y=224440
X858 1632 1266 11 10 37 482 MXI2XL $T=227940 209380 0 0 $X=227340 $Y=209020
X859 1633 1265 11 10 39 479 MXI2XL $T=233160 292900 0 180 $X=227920 $Y=287080
X860 475 1259 11 10 37 1634 MXI2XL $T=230840 240700 1 0 $X=230240 $Y=234880
X861 1591 1262 11 10 39 1635 MXI2XL $T=233740 272020 1 0 $X=233140 $Y=266200
X862 486 1267 11 10 39 494 MXI2XL $T=240120 282460 0 180 $X=234880 $Y=276640
X863 488 1269 11 10 37 1450 MXI2XL $T=246500 230260 0 0 $X=245900 $Y=229900
X864 1636 1275 11 10 37 490 MXI2XL $T=262160 230260 1 180 $X=256920 $Y=229900
X865 493 1274 11 10 37 496 MXI2XL $T=263900 230260 0 0 $X=263300 $Y=229900
X866 1637 1273 11 10 39 1638 MXI2XL $T=268540 272020 0 0 $X=267940 $Y=271660
X867 1639 1279 11 10 39 1640 MXI2XL $T=281300 324220 0 180 $X=276060 $Y=318400
X868 1451 1277 11 10 168 501 MXI2XL $T=277820 209380 0 0 $X=277220 $Y=209020
X869 491 1276 11 10 168 498 MXI2XL $T=278400 198940 1 0 $X=277800 $Y=193120
X870 1453 1282 11 10 190 521 MXI2XL $T=316680 272020 0 180 $X=311440 $Y=266200
X871 527 1283 11 10 190 1641 MXI2XL $T=329440 261580 1 0 $X=328840 $Y=255760
X872 1642 1284 11 10 190 529 MXI2XL $T=335820 240700 1 180 $X=330580 $Y=240340
X873 194 1285 11 10 168 532 MXI2XL $T=332920 209380 1 0 $X=332320 $Y=203560
X874 535 1287 11 10 198 534 MXI2XL $T=338140 365980 0 180 $X=332900 $Y=360160
X875 1643 1288 11 10 199 1644 MXI2XL $T=341040 313780 0 180 $X=335800 $Y=307960
X876 1600 1292 11 10 198 1645 MXI2XL $T=346840 365980 0 180 $X=341600 $Y=360160
X877 542 1290 11 10 199 530 MXI2XL $T=352060 313780 0 180 $X=346820 $Y=307960
X878 1646 1289 11 10 198 553 MXI2XL $T=353800 334660 0 0 $X=353200 $Y=334300
X879 556 1294 11 10 190 557 MXI2XL $T=360180 209380 1 180 $X=354940 $Y=209020
X880 1462 1295 11 10 199 560 MXI2XL $T=356120 313780 1 0 $X=355520 $Y=307960
X881 1647 1296 11 10 199 1648 MXI2XL $T=370040 282460 0 180 $X=364800 $Y=276640
X882 1649 1299 11 10 190 1650 MXI2XL $T=385700 209380 0 180 $X=380460 $Y=203560
X883 1604 1305 11 10 190 1651 MXI2XL $T=394980 209380 0 180 $X=389740 $Y=203560
X884 586 1311 11 10 190 581 MXI2XL $T=408320 240700 1 0 $X=407720 $Y=234880
X885 624 1307 11 10 198 1375 MXI2XL $T=418760 345100 0 180 $X=413520 $Y=339280
X886 235 1315 11 10 190 236 MXI2XL $T=422240 209380 1 180 $X=417000 $Y=209020
X887 644 1316 11 10 199 632 MXI2XL $T=438480 261580 0 180 $X=433240 $Y=255760
X888 1652 1323 11 10 190 1489 MXI2XL $T=445440 198940 0 0 $X=444840 $Y=198580
X889 1383 1327 11 10 199 689 MXI2XL $T=459940 272020 1 180 $X=454700 $Y=271660
X890 1653 282 11 10 283 284 MXI2XL $T=488940 365980 0 0 $X=488340 $Y=365620
X891 1381 1335 11 10 198 1581 MXI2XL $T=494740 345100 1 180 $X=489500 $Y=344740
X892 1654 1337 11 10 198 1655 MXI2XL $T=506340 292900 0 180 $X=501100 $Y=287080
X893 1656 1342 11 10 199 301 MXI2XL $T=526060 219820 1 180 $X=520820 $Y=219460
X894 1657 1341 11 10 199 1658 MXI2XL $T=527800 219820 0 180 $X=522560 $Y=214000
X895 1659 1344 11 10 198 1660 MXI2XL $T=527800 324220 1 180 $X=522560 $Y=323860
X896 1661 1475 11 10 1480 631 AND3X1 $T=410060 272020 0 0 $X=409460 $Y=271660
X897 1619 11 10 1415 1108 1662 783 37 AOI221XL $T=89320 230260 1 180 $X=82920 $Y=229900
X898 1587 11 10 1425 1109 1663 818 1538 AOI221XL $T=139200 219820 1 0 $X=138600 $Y=214000
X899 1111 11 10 1143 387 1664 1426 39 AOI221XL $T=146740 282460 1 180 $X=140340 $Y=282100
X900 1665 11 10 1428 1112 1408 1173 1666 AOI221XL $T=160660 282460 1 180 $X=154260 $Y=282100
X901 1667 11 10 1432 1177 1406 1101 1544 AOI221XL $T=169940 261580 0 180 $X=163540 $Y=255760
X902 1124 11 10 821 1668 1669 1433 1546 AOI221XL $T=178640 209380 0 0 $X=178040 $Y=209020
X903 1176 11 10 1118 432 1670 1436 98 AOI221XL $T=188500 272020 0 0 $X=187900 $Y=271660
X904 1123 11 10 848 482 1671 1447 54 AOI221XL $T=239540 219820 0 180 $X=233140 $Y=214000
X905 175 11 10 898 194 1672 1455 168 AOI221XL $T=325960 209380 1 0 $X=325360 $Y=203560
X906 1600 11 10 1460 1286 1673 925 198 AOI221XL $T=352640 345100 0 0 $X=352040 $Y=344740
X907 1647 11 10 1461 1213 1674 934 199 AOI221XL $T=365400 282460 0 180 $X=359000 $Y=276640
X908 208 11 10 963 586 1675 1478 190 AOI221XL $T=408320 240700 0 180 $X=401920 $Y=234880
X909 206 11 10 955 1676 581 1491 1569 AOI221XL $T=413540 230260 1 0 $X=412940 $Y=224440
X910 1605 11 10 1493 227 1652 232 1570 AOI221XL $T=424560 198940 1 180 $X=418160 $Y=198580
X911 1317 11 10 986 1375 1677 1494 222 AOI221XL $T=420500 324220 0 0 $X=419900 $Y=323860
X912 632 11 10 1492 1212 1678 994 231 AOI221XL $T=430940 261580 0 180 $X=424540 $Y=255760
X913 219 11 10 992 1489 1679 1495 209 AOI221XL $T=439640 198940 1 180 $X=433240 $Y=198580
X914 1383 11 10 1503 1210 1680 1000 199 AOI221XL $T=452400 282460 1 0 $X=451800 $Y=276640
X915 1328 11 10 1027 1381 1681 1509 198 AOI221XL $T=484880 345100 1 0 $X=484280 $Y=339280
X916 1328 11 10 1063 1659 1682 1531 198 AOI221XL $T=518520 313780 0 0 $X=517920 $Y=313420
X917 1384 353 11 10 354 1683 54 62 BMXIX2 $T=91060 198940 0 0 $X=90460 $Y=198580
X918 1684 367 11 10 368 1685 39 789 BMXIX2 $T=106140 272020 1 180 $X=90460 $Y=271660
X919 1686 447 11 10 448 1687 39 837 BMXIX2 $T=203580 261580 0 0 $X=202980 $Y=261220
X920 1688 502 11 10 503 1561 186 905 BMXIX2 $T=293480 230260 1 0 $X=292880 $Y=224440
X921 1371 178 11 10 507 1689 186 890 BMXIX2 $T=297540 209380 1 0 $X=296940 $Y=203560
X922 1392 514 11 10 515 1690 186 887 BMXIX2 $T=308560 219820 1 0 $X=307960 $Y=214000
X923 1373 537 11 10 538 1691 209 921 BMXIX2 $T=342200 261580 0 0 $X=341600 $Y=261220
X924 1692 547 11 10 548 1564 209 944 BMXIX2 $T=359020 261580 0 0 $X=358420 $Y=261220
X925 1393 551 11 10 552 1693 209 941 BMXIX2 $T=360760 261580 1 0 $X=360160 $Y=255760
X926 1396 621 11 10 622 1694 231 1007 BMXIX2 $T=415860 292900 0 0 $X=415260 $Y=292540
X927 1377 627 11 10 628 1695 222 246 BMXIX2 $T=425140 365980 0 0 $X=424540 $Y=365620
X928 1696 653 11 10 654 1398 222 239 BMXIX2 $T=449500 313780 0 180 $X=433820 $Y=307960
X929 1697 655 11 10 656 1573 222 248 BMXIX2 $T=454140 365980 0 180 $X=438460 $Y=360160
X930 1576 694 11 10 695 1698 222 243 BMXIX2 $T=465160 334660 0 180 $X=449480 $Y=328840
X931 1399 684 11 10 685 1699 199 1017 BMXIX2 $T=450660 261580 1 0 $X=450060 $Y=255760
X932 1401 677 11 10 678 1700 222 263 BMXIX2 $T=450660 365980 0 0 $X=450060 $Y=365620
X933 1575 269 11 10 715 267 209 1034 BMXIX2 $T=468060 188500 0 0 $X=467460 $Y=188140
X934 1402 270 11 10 710 1701 190 1022 BMXIX2 $T=468060 198940 0 0 $X=467460 $Y=198580
X935 1702 724 11 10 725 1379 222 265 BMXIX2 $T=483140 334660 0 180 $X=467460 $Y=328840
X936 1582 787 11 10 1109 353 ADDHX1 $T=108460 209380 0 0 $X=107860 $Y=209020
X937 1703 812 11 10 1112 367 ADDHX1 $T=109040 282460 0 0 $X=108440 $Y=282100
X938 1403 806 11 10 1108 70 ADDHX1 $T=126440 219820 0 180 $X=116560 $Y=214000
X939 1420 808 11 10 1109 379 ADDHX1 $T=120060 209380 1 0 $X=119460 $Y=203560
X940 1704 1116 11 10 91 1705 ADDHX1 $T=151960 345100 0 180 $X=142080 $Y=339280
X941 1706 91 11 10 1115 1707 ADDHX1 $T=143840 355540 1 0 $X=143240 $Y=349720
X942 1708 1141 11 10 91 1709 ADDHX1 $T=186180 345100 1 180 $X=176300 $Y=344740
X943 1710 1141 11 10 83 1711 ADDHX1 $T=182120 334660 1 0 $X=181520 $Y=328840
X944 1439 826 11 10 1124 119 ADDHX1 $T=186760 188500 0 0 $X=186160 $Y=188140
X945 437 830 11 10 1123 123 ADDHX1 $T=198360 188500 0 0 $X=197760 $Y=188140
X946 1712 1133 11 10 1176 447 ADDHX1 $T=198360 282460 1 0 $X=197760 $Y=276640
X947 455 131 11 10 1152 461 ADDHX1 $T=210540 334660 1 0 $X=209940 $Y=328840
X948 1593 835 11 10 1124 127 ADDHX1 $T=211120 198940 1 0 $X=210520 $Y=193120
X949 1713 141 11 10 121 766 ADDHX1 $T=229100 365980 1 180 $X=219220 $Y=365620
X950 1714 131 11 10 1153 1715 ADDHX1 $T=220980 334660 0 0 $X=220380 $Y=334300
X951 1716 143 11 10 1153 1717 ADDHX1 $T=239540 313780 1 180 $X=229660 $Y=313420
X952 1370 174 11 10 175 502 ADDHX1 $T=297540 209380 0 180 $X=287660 $Y=203560
X953 505 853 11 10 182 514 ADDHX1 $T=297540 219820 1 0 $X=296940 $Y=214000
X954 1457 888 11 10 206 537 ADDHX1 $T=353800 240700 1 180 $X=343920 $Y=240340
X955 1372 904 11 10 208 547 ADDHX1 $T=349740 261580 1 0 $X=349140 $Y=255760
X956 1718 885 11 10 206 551 ADDHX1 $T=366560 251140 0 0 $X=365960 $Y=250780
X957 1476 919 11 10 1211 579 ADDHX1 $T=385120 313780 0 0 $X=384520 $Y=313420
X958 1409 943 11 10 1210 607 ADDHX1 $T=401360 313780 0 0 $X=400760 $Y=313420
X959 1608 939 11 10 1211 621 ADDHX1 $T=421080 313780 1 0 $X=420480 $Y=307960
X960 1497 1208 11 10 1312 627 ADDHX1 $T=436160 355540 1 180 $X=426280 $Y=355180
X961 1376 1207 11 10 1328 655 ADDHX1 $T=436160 355540 1 0 $X=435560 $Y=349720
X962 670 1005 11 10 1312 677 ADDHX1 $T=444280 376420 1 0 $X=443680 $Y=370600
X963 686 1015 11 10 1286 653 ADDHX1 $T=460520 313780 0 180 $X=450640 $Y=307960
X964 1612 1020 11 10 1213 684 ADDHX1 $T=465740 251140 0 180 $X=455860 $Y=245320
X965 1378 1216 11 10 1317 694 ADDHX1 $T=477340 324220 1 180 $X=467460 $Y=323860
X966 1411 274 11 10 1212 706 ADDHX1 $T=482560 251140 1 180 $X=472680 $Y=250780
X967 1516 1218 11 10 1286 724 ADDHX1 $T=486620 334660 1 0 $X=486020 $Y=328840
X968 1514 279 11 10 1213 732 ADDHX1 $T=487200 251140 1 0 $X=486600 $Y=245320
X969 37 11 10 1719 1662 1227 AO21X1 $T=89320 240700 0 180 $X=83500 $Y=234880
X970 357 11 10 1720 54 1721 AO21X1 $T=97440 219820 0 180 $X=91620 $Y=214000
X971 1108 11 10 1413 1620 1720 AO21X1 $T=92220 230260 1 0 $X=91620 $Y=224440
X972 1109 11 10 793 355 1385 AO21X1 $T=95700 209380 1 0 $X=95100 $Y=203560
X973 1109 11 10 361 358 388 AO21X1 $T=100920 219820 0 0 $X=100320 $Y=219460
X974 1111 11 10 374 364 1722 AO21X1 $T=113680 292900 1 180 $X=107860 $Y=292540
X975 1109 11 10 372 1385 377 AO21X1 $T=110200 209380 1 0 $X=109600 $Y=203560
X976 39 11 10 1723 1664 1242 AO21X1 $T=143840 282460 0 180 $X=138020 $Y=276640
X977 389 11 10 1663 54 1724 AO21X1 $T=139780 209380 0 0 $X=139180 $Y=209020
X978 404 11 10 1725 98 1726 AO21X1 $T=156600 272020 0 180 $X=150780 $Y=266200
X979 1122 11 10 1116 91 1543 AO21X1 $T=153700 355540 1 0 $X=153100 $Y=349720
X980 1112 11 10 409 386 1727 AO21X1 $T=160080 292900 1 0 $X=159480 $Y=287080
X981 407 11 10 1727 39 1728 AO21X1 $T=162400 282460 0 0 $X=161800 $Y=282100
X982 454 11 10 1669 37 1729 AO21X1 $T=180960 209380 0 180 $X=175140 $Y=203560
X983 1151 11 10 1141 91 1730 AO21X1 $T=185020 355540 1 0 $X=184420 $Y=349720
X984 1151 11 10 1141 83 1731 AO21X1 $T=191400 334660 1 180 $X=185580 $Y=334300
X985 98 11 10 1732 1670 1255 AO21X1 $T=190820 261580 0 0 $X=190220 $Y=261220
X986 1177 11 10 428 431 1725 AO21X1 $T=190820 272020 1 0 $X=190220 $Y=266200
X987 1124 11 10 1441 1391 1438 AO21X1 $T=210540 198940 1 180 $X=204720 $Y=198580
X988 1123 11 10 1441 463 1387 AO21X1 $T=211120 209380 0 180 $X=205300 $Y=203560
X989 1123 11 10 1445 468 443 AO21X1 $T=215760 198940 1 180 $X=209940 $Y=198580
X990 1124 11 10 1445 466 453 AO21X1 $T=218080 209380 0 180 $X=212260 $Y=203560
X991 1167 11 10 131 1153 1733 AO21X1 $T=220980 345100 1 180 $X=215160 $Y=344740
X992 1124 11 10 1448 481 473 AO21X1 $T=225040 219820 0 180 $X=219220 $Y=214000
X993 1177 11 10 460 1635 1734 AO21X1 $T=219820 282460 1 0 $X=219220 $Y=276640
X994 1124 11 10 844 473 1391 AO21X1 $T=226200 198940 1 180 $X=220380 $Y=198580
X995 844 11 10 1123 1735 463 AO21X1 $T=227940 209380 1 180 $X=222120 $Y=209020
X996 465 11 10 1735 37 1736 AO21X1 $T=224460 209380 1 0 $X=223860 $Y=203560
X997 1123 11 10 1448 1632 1735 AO21X1 $T=230840 219820 0 180 $X=225020 $Y=214000
X998 54 11 10 1737 1671 1268 AO21X1 $T=240700 209380 1 0 $X=240100 $Y=203560
X999 1193 11 10 143 1153 1555 AO21X1 $T=245920 334660 0 180 $X=240100 $Y=328840
X1000 163 11 10 1192 1153 1560 AO21X1 $T=257520 334660 0 0 $X=256920 $Y=334300
X1001 506 11 10 512 179 1688 AO21X1 $T=294640 209380 1 180 $X=288820 $Y=209020
X1002 175 11 10 1452 509 181 AO21X1 $T=290000 198940 1 0 $X=289400 $Y=193120
X1003 853 11 10 175 509 1562 AO21X1 $T=290000 198940 0 0 $X=289400 $Y=198580
X1004 182 11 10 1452 513 510 AO21X1 $T=297540 188500 0 0 $X=296940 $Y=188140
X1005 182 11 10 516 519 183 AO21X1 $T=301600 198940 1 0 $X=301000 $Y=193120
X1006 518 11 10 525 186 1738 AO21X1 $T=317840 198940 1 180 $X=312020 $Y=198580
X1007 168 11 10 1739 1672 1291 AO21X1 $T=339880 209380 1 0 $X=339280 $Y=203560
X1008 206 11 10 1456 1395 539 AO21X1 $T=352640 251140 0 180 $X=346820 $Y=245320
X1009 208 11 10 1456 566 549 AO21X1 $T=353220 251140 1 0 $X=352620 $Y=245320
X1010 888 11 10 208 549 1346 AO21X1 $T=354960 240700 0 0 $X=354360 $Y=240340
X1011 198 11 10 1740 1673 1293 AO21X1 $T=360180 355540 1 180 $X=354360 $Y=355180
X1012 885 11 10 208 566 1565 AO21X1 $T=364240 251140 1 0 $X=363640 $Y=245320
X1013 206 11 10 894 1741 1395 AO21X1 $T=365980 240700 0 0 $X=365380 $Y=240340
X1014 199 11 10 1742 1674 1301 AO21X1 $T=370040 282460 1 0 $X=369440 $Y=276640
X1015 1286 11 10 564 1645 1743 AO21X1 $T=370620 355540 0 0 $X=370020 $Y=355180
X1016 1394 11 10 1741 190 1744 AO21X1 $T=378160 240700 1 0 $X=377560 $Y=234880
X1017 597 11 10 1743 222 1745 AO21X1 $T=389180 355540 1 180 $X=383360 $Y=355180
X1018 1213 11 10 1467 1648 1746 AO21X1 $T=392660 272020 1 180 $X=386840 $Y=271660
X1019 951 11 10 1286 1743 1747 AO21X1 $T=389180 355540 0 0 $X=388580 $Y=355180
X1020 206 11 10 575 585 1741 AO21X1 $T=393820 240700 1 0 $X=393220 $Y=234880
X1021 957 11 10 227 1651 1748 AO21X1 $T=400200 209380 0 180 $X=394380 $Y=203560
X1022 968 11 10 1212 577 1354 AO21X1 $T=404840 261580 1 180 $X=399020 $Y=261220
X1023 588 11 10 1749 231 1750 AO21X1 $T=399620 303340 0 0 $X=399020 $Y=302980
X1024 1479 11 10 1751 190 1752 AO21X1 $T=400200 230260 1 0 $X=399600 $Y=224440
X1025 1475 11 10 1746 231 1753 AO21X1 $T=406000 282460 0 180 $X=400180 $Y=276640
X1026 968 11 10 1213 1746 615 AO21X1 $T=406580 272020 1 180 $X=400760 $Y=271660
X1027 1211 11 10 610 1397 605 AO21X1 $T=414120 313780 0 180 $X=408300 $Y=307960
X1028 612 11 10 1748 209 1754 AO21X1 $T=410640 198940 1 0 $X=410040 $Y=193120
X1029 190 11 10 1755 1675 1309 AO21X1 $T=418180 240700 0 180 $X=412360 $Y=234880
X1030 1210 11 10 1483 636 593 AO21X1 $T=421080 292900 0 180 $X=415260 $Y=287080
X1031 1211 11 10 1483 640 587 AO21X1 $T=422240 303340 0 180 $X=416420 $Y=297520
X1032 222 11 10 1756 1677 1318 AO21X1 $T=425720 334660 0 180 $X=419900 $Y=328840
X1033 1211 11 10 979 633 1397 AO21X1 $T=429780 282460 1 180 $X=423960 $Y=282100
X1034 1208 11 10 1328 637 1356 AO21X1 $T=433260 345100 1 180 $X=427440 $Y=344740
X1035 231 11 10 1757 1678 1319 AO21X1 $T=430360 251140 0 0 $X=429760 $Y=250780
X1036 1328 11 10 1500 676 637 AO21X1 $T=443700 345100 1 180 $X=437880 $Y=344740
X1037 639 11 10 646 231 1758 AO21X1 $T=439060 292900 0 0 $X=438460 $Y=292540
X1038 209 11 10 1759 1679 1321 AO21X1 $T=440220 198940 0 0 $X=439620 $Y=198580
X1039 1312 11 10 1500 669 641 AO21X1 $T=445440 355540 1 180 $X=439620 $Y=355180
X1040 1213 11 10 648 631 663 AO21X1 $T=440800 261580 1 0 $X=440200 $Y=255760
X1041 1005 11 10 1328 676 1574 AO21X1 $T=444860 345100 0 0 $X=444260 $Y=344740
X1042 659 11 10 662 198 1760 AO21X1 $T=450660 324220 1 180 $X=444840 $Y=323860
X1043 682 11 10 652 199 1761 AO21X1 $T=446020 251140 1 0 $X=445420 $Y=245320
X1044 1328 11 10 1504 703 617 AO21X1 $T=448340 355540 0 0 $X=447740 $Y=355180
X1045 1312 11 10 1504 699 625 AO21X1 $T=448920 355540 1 0 $X=448320 $Y=349720
X1046 254 11 10 667 190 1762 AO21X1 $T=452400 198940 0 0 $X=451800 $Y=198580
X1047 1213 11 10 1008 663 1400 AO21X1 $T=452400 251140 0 0 $X=451800 $Y=250780
X1048 1317 11 10 672 650 728 AO21X1 $T=453560 324220 1 0 $X=452960 $Y=318400
X1049 671 11 10 668 617 1697 AO21X1 $T=454140 365980 1 0 $X=453540 $Y=360160
X1050 687 11 10 692 728 1698 AO21X1 $T=461100 324220 1 180 $X=455280 $Y=323860
X1051 199 11 10 1763 1680 1325 AO21X1 $T=458200 282460 1 0 $X=457600 $Y=276640
X1052 1212 11 10 1505 680 716 AO21X1 $T=460520 240700 1 0 $X=459920 $Y=234880
X1053 1213 11 10 1505 683 718 AO21X1 $T=460520 240700 0 0 $X=459920 $Y=240340
X1054 1015 11 10 1317 697 1577 AO21X1 $T=460520 313780 1 0 $X=459920 $Y=307960
X1055 1317 11 10 1508 697 704 AO21X1 $T=468060 313780 1 0 $X=467460 $Y=307960
X1056 1286 11 10 1508 693 722 AO21X1 $T=468060 324220 1 0 $X=467460 $Y=318400
X1057 698 11 10 1764 222 1765 AO21X1 $T=468060 355540 1 0 $X=467460 $Y=349720
X1058 1213 11 10 714 1400 720 AO21X1 $T=473280 251140 1 0 $X=472680 $Y=245320
X1059 1218 11 10 1317 704 1361 AO21X1 $T=478500 313780 0 180 $X=472680 $Y=307960
X1060 719 11 10 1766 199 1767 AO21X1 $T=485460 230260 1 180 $X=479640 $Y=229900
X1061 1328 11 10 727 1581 1764 AO21X1 $T=484880 345100 0 0 $X=484280 $Y=344740
X1062 198 11 10 1768 1681 1331 AO21X1 $T=497640 345100 0 180 $X=491820 $Y=339280
X1063 286 11 10 245 1653 291 AO21X1 $T=497640 376420 1 0 $X=497040 $Y=370600
X1064 1046 11 10 1328 750 1364 AO21X1 $T=498220 324220 1 0 $X=497620 $Y=318400
X1065 1046 11 10 1312 1769 1770 AO21X1 $T=502860 324220 0 0 $X=502260 $Y=323860
X1066 1049 11 10 1210 738 1368 AO21X1 $T=512140 230260 1 180 $X=506320 $Y=229900
X1067 742 11 10 1769 198 1771 AO21X1 $T=513880 324220 1 180 $X=508060 $Y=323860
X1068 1210 11 10 1527 301 738 AO21X1 $T=509820 219820 0 0 $X=509220 $Y=219460
X1069 752 11 10 1772 199 1773 AO21X1 $T=519680 240700 1 180 $X=513860 $Y=240340
X1070 1049 11 10 1211 1772 1774 AO21X1 $T=517940 240700 1 0 $X=517340 $Y=234880
X1071 1328 11 10 1526 1660 750 AO21X1 $T=517940 324220 0 0 $X=517340 $Y=323860
X1072 198 11 10 1775 1682 1345 AO21X1 $T=527800 324220 0 0 $X=527200 $Y=323860
X1073 786 800 11 10 796 XNOR2X1 $T=93380 240700 1 0 $X=92780 $Y=234880
X1074 801 1126 11 10 1085 XNOR2X1 $T=117160 355540 0 180 $X=110180 $Y=349720
X1075 1110 1111 11 10 1177 XNOR2X1 $T=152540 261580 0 180 $X=145560 $Y=255760
X1076 1107 1707 11 10 1776 XNOR2X1 $T=156020 345100 1 180 $X=149040 $Y=344740
X1077 1106 1705 11 10 1588 XNOR2X1 $T=151960 345100 1 0 $X=151360 $Y=339280
X1078 108 1123 11 10 1109 XNOR2X1 $T=171680 209380 0 180 $X=164700 $Y=203560
X1079 1135 1711 11 10 1589 XNOR2X1 $T=189080 324220 1 180 $X=182100 $Y=323860
X1080 1134 1709 11 10 1590 XNOR2X1 $T=183860 345100 1 0 $X=183260 $Y=339280
X1081 1161 1717 11 10 1597 XNOR2X1 $T=230260 313780 1 180 $X=223280 $Y=313420
X1082 852 765 11 10 1162 XNOR2X1 $T=233160 292900 1 0 $X=232560 $Y=287080
X1083 154 851 11 10 856 XNOR2X1 $T=244180 240700 0 0 $X=243580 $Y=240340
X1084 881 842 11 10 854 XNOR2X1 $T=276660 209380 1 180 $X=269680 $Y=209020
X1085 918 880 11 10 894 XNOR2X1 $T=338140 261580 1 0 $X=337540 $Y=255760
X1086 947 917 11 10 939 XNOR2X1 $T=375840 313780 0 180 $X=368860 $Y=307960
X1087 225 1207 11 10 945 XNOR2X1 $T=390340 345100 1 180 $X=383360 $Y=344740
X1088 629 206 11 10 227 XNOR2X1 $T=424560 209380 0 0 $X=423960 $Y=209020
X1089 251 1312 11 10 1286 XNOR2X1 $T=447180 365980 1 180 $X=440200 $Y=365620
X1090 690 1210 11 10 1213 XNOR2X1 $T=447760 282460 1 180 $X=440780 $Y=282100
X1091 762 1021 11 10 1018 XNOR2X1 $T=475600 219820 1 180 $X=468620 $Y=219460
X1092 259 761 11 10 1215 XNOR2X1 $T=471540 303340 1 0 $X=470940 $Y=297520
X1093 37 11 10 352 356 1721 1230 OAI31XL $T=89320 209380 1 180 $X=84080 $Y=209020
X1094 385 11 10 376 1777 1724 94 OAI31XL $T=139200 209380 1 0 $X=138600 $Y=203560
X1095 98 11 10 1666 1665 1728 1246 OAI31XL $T=167040 282460 0 180 $X=161800 $Y=276640
X1096 39 11 10 1544 1667 1726 1247 OAI31XL $T=172260 261580 1 180 $X=167020 $Y=261220
X1097 423 11 10 440 1778 1729 414 OAI31XL $T=180380 198940 1 180 $X=175140 $Y=198580
X1098 54 11 10 468 474 1736 1263 OAI31XL $T=229680 198940 0 0 $X=229080 $Y=198580
X1099 168 11 10 522 1599 1738 1281 OAI31XL $T=317260 209380 0 180 $X=312020 $Y=203560
X1100 544 11 10 545 1779 209 1780 OAI31XL $T=360180 230260 0 0 $X=359580 $Y=229900
X1101 209 11 10 562 1347 1780 1214 OAI31XL $T=374680 230260 1 180 $X=369440 $Y=229900
X1102 209 11 10 570 1602 1744 1300 OAI31XL $T=379320 240700 0 0 $X=378720 $Y=240340
X1103 198 11 10 572 1601 1745 1302 OAI31XL $T=379320 355540 0 0 $X=378720 $Y=355180
X1104 199 11 10 584 578 1753 1304 OAI31XL $T=395560 282460 1 0 $X=394960 $Y=276640
X1105 590 11 10 604 1781 1750 1782 OAI31XL $T=402520 292900 0 0 $X=401920 $Y=292540
X1106 209 11 10 1569 1676 1752 1314 OAI31XL $T=406580 230260 1 0 $X=405980 $Y=224440
X1107 190 11 10 1570 1605 1754 1310 OAI31XL $T=417020 198940 1 180 $X=411780 $Y=198580
X1108 619 11 10 617 1783 222 1784 OAI31XL $T=418180 365980 1 0 $X=417580 $Y=360160
X1109 222 11 10 625 1357 1784 241 OAI31XL $T=424560 365980 1 0 $X=423960 $Y=360160
X1110 199 11 10 636 634 1758 1320 OAI31XL $T=430940 292900 0 0 $X=430340 $Y=292540
X1111 222 11 10 650 1609 1760 1322 OAI31XL $T=439060 324220 0 0 $X=438460 $Y=323860
X1112 231 11 10 680 664 1761 1324 OAI31XL $T=447180 251140 0 0 $X=446580 $Y=250780
X1113 209 11 10 255 1611 1762 1326 OAI31XL $T=453560 198940 1 0 $X=452960 $Y=193120
X1114 712 11 10 709 1785 1767 1786 OAI31XL $T=474440 230260 1 180 $X=469200 $Y=229900
X1115 198 11 10 703 1613 1765 1329 OAI31XL $T=469800 355540 0 0 $X=469200 $Y=355180
X1116 198 11 10 701 1362 1787 273 OAI31XL $T=483140 324220 0 180 $X=477900 $Y=318400
X1117 734 11 10 728 1788 198 1787 OAI31XL $T=489520 324220 0 180 $X=484280 $Y=318400
X1118 231 11 10 745 739 1773 1336 OAI31XL $T=498800 240700 1 0 $X=498200 $Y=234880
X1119 222 11 10 749 751 1771 1340 OAI31XL $T=512140 334660 1 0 $X=511540 $Y=328840
X1120 1534 384 11 10 1421 37 1424 AOI31XL $T=129340 209380 1 0 $X=128740 $Y=203560
X1121 444 422 11 10 1440 54 1435 AOI31XL $T=192560 198940 1 180 $X=187320 $Y=198580
X1122 546 543 11 10 1458 190 1463 AOI31XL $T=347420 230260 0 0 $X=346820 $Y=229900
X1123 594 589 11 10 1477 199 1472 AOI31XL $T=398460 292900 1 180 $X=393220 $Y=292540
X1124 597 600 11 10 1747 222 1474 AOI31XL $T=402520 355540 1 180 $X=397280 $Y=355180
X1125 1475 1480 11 10 615 231 1482 AOI31XL $T=406580 282460 1 0 $X=405980 $Y=276640
X1126 618 620 11 10 1498 198 1486 AOI31XL $T=417020 355540 1 180 $X=411780 $Y=355180
X1127 717 711 11 10 1515 231 1521 AOI31XL $T=487780 240700 1 0 $X=487180 $Y=234880
X1128 729 735 11 10 1517 222 1518 AOI31XL $T=493580 324220 1 180 $X=488340 $Y=323860
X1129 742 747 11 10 1770 198 1525 AOI31XL $T=516780 345100 0 180 $X=511540 $Y=339280
X1130 752 755 11 10 1774 199 1529 AOI31XL $T=524320 251140 0 180 $X=519080 $Y=245320
X1131 794 1109 11 10 1683 358 1584 AOI211XL $T=96860 219820 0 0 $X=96260 $Y=219460
X1132 812 1111 11 10 386 1535 1586 AOI211XL $T=126440 292900 1 180 $X=121780 $Y=292540
X1133 806 1109 11 10 1404 388 1585 AOI211XL $T=126440 219820 1 0 $X=125840 $Y=214000
X1134 1430 1541 11 10 1249 1540 1789 AOI211XL $T=157760 334660 1 0 $X=157160 $Y=328840
X1135 1731 435 11 10 1250 1710 426 AOI211XL $T=184440 334660 1 180 $X=179780 $Y=334300
X1136 1730 441 11 10 1542 1708 430 AOI211XL $T=187920 345100 0 0 $X=187320 $Y=344740
X1137 1133 1177 11 10 1631 1550 1592 AOI211XL $T=200680 272020 0 0 $X=200080 $Y=271660
X1138 1733 449 11 10 1261 1714 458 AOI211XL $T=211120 345100 1 0 $X=210520 $Y=339280
X1139 845 1124 11 10 125 466 464 AOI211XL $T=218080 209380 1 0 $X=217480 $Y=203560
X1140 1449 1554 11 10 1270 1556 1790 AOI211XL $T=245920 324220 0 0 $X=245320 $Y=323860
X1141 174 182 11 10 1689 183 504 AOI211XL $T=295800 198940 1 0 $X=295200 $Y=193120
X1142 863 182 11 10 1690 519 508 AOI211XL $T=310880 198940 0 180 $X=306220 $Y=193120
X1143 904 206 11 10 1691 562 550 AOI211XL $T=352640 251140 0 0 $X=352040 $Y=250780
X1144 895 206 11 10 1693 570 565 AOI211XL $T=371780 251140 1 0 $X=371180 $Y=245320
X1145 943 1211 11 10 1410 587 1603 AOI211XL $T=401360 303340 1 0 $X=400760 $Y=297520
X1146 980 1211 11 10 1694 640 1606 AOI211XL $T=422820 303340 1 0 $X=422220 $Y=297520
X1147 1207 1312 11 10 1695 625 638 AOI211XL $T=431520 355540 1 0 $X=430920 $Y=349720
X1148 1012 1286 11 10 1696 660 696 AOI211XL $T=450080 313780 0 0 $X=449480 $Y=313420
X1149 1009 1213 11 10 1699 683 1610 AOI211XL $T=454140 240700 0 0 $X=453540 $Y=240340
X1150 1003 1312 11 10 1700 699 675 AOI211XL $T=455300 355540 1 0 $X=454700 $Y=349720
X1151 250 227 11 10 1701 665 681 AOI211XL $T=457620 198940 0 0 $X=457020 $Y=198580
X1152 1216 1286 11 10 1702 701 705 AOI211XL $T=477340 324220 0 180 $X=472680 $Y=318400
X1153 274 1213 11 10 1412 718 1615 AOI211XL $T=484880 240700 1 180 $X=480220 $Y=240340
X1154 439 11 10 438 1438 122 1386 54 AOI32XL $T=200100 198940 1 0 $X=199500 $Y=193120
X1155 774 11 10 30 43 339 ACHCONX2 $T=44660 198940 1 0 $X=44080 $Y=193120
X1156 783 11 10 778 1616 335 ACHCONX2 $T=46980 230260 1 0 $X=46400 $Y=224440
X1157 757 11 10 768 341 1616 ACHCONX2 $T=46980 261580 1 0 $X=46400 $Y=255760
X1158 794 11 10 771 1624 341 ACHCONX2 $T=48140 261580 0 0 $X=47560 $Y=261220
X1159 757 11 10 769 345 333 ACHCONX2 $T=48140 272020 1 0 $X=47560 $Y=266200
X1160 25 11 10 1093 343 338 ACHCONX2 $T=48140 345100 1 0 $X=47560 $Y=339280
X1161 782 11 10 778 333 1417 ACHCONX2 $T=48720 240700 1 0 $X=48140 $Y=234880
X1162 1072 11 10 1078 369 344 ACHCONX2 $T=56260 324220 0 0 $X=55680 $Y=323860
X1163 1093 11 10 1100 1618 1621 ACHCONX2 $T=56840 313780 0 0 $X=56260 $Y=313420
X1164 772 11 10 794 1623 346 ACHCONX2 $T=58000 272020 0 0 $X=57420 $Y=271660
X1165 1077 11 10 1112 359 1618 ACHCONX2 $T=87000 292900 1 180 $X=57420 $Y=292540
X1166 1075 11 10 1082 337 1533 ACHCONX2 $T=98020 355540 0 180 $X=68440 $Y=349720
X1167 1108 11 10 782 1719 1620 ACHCONX2 $T=70180 240700 0 0 $X=69600 $Y=240340
X1168 1092 11 10 1100 349 1622 ACHCONX2 $T=72500 313780 1 0 $X=71920 $Y=307960
X1169 26 11 10 41 339 1416 ACHCONX2 $T=73660 198940 1 0 $X=73080 $Y=193120
X1170 1073 11 10 1078 365 347 ACHCONX2 $T=75980 334660 0 0 $X=75400 $Y=334300
X1171 1076 11 10 1082 1617 1532 ACHCONX2 $T=76560 355540 0 0 $X=75980 $Y=355180
X1172 787 11 10 790 1791 1623 ACHCONX2 $T=77140 261580 1 0 $X=76560 $Y=255760
X1173 787 11 10 791 1792 1624 ACHCONX2 $T=77140 261580 0 0 $X=76560 $Y=261220
X1174 1111 11 10 1097 1685 359 ACHCONX2 $T=77140 292900 1 0 $X=76560 $Y=287080
X1175 1111 11 10 1077 363 350 ACHCONX2 $T=77140 303340 1 0 $X=76560 $Y=297520
X1176 1111 11 10 1096 1684 364 ACHCONX2 $T=77140 303340 0 0 $X=76560 $Y=302980
X1177 1088 11 10 1097 380 370 ACHCONX2 $T=77140 324220 1 0 $X=76560 $Y=318400
X1178 1092 11 10 25 347 1617 ACHCONX2 $T=77140 345100 1 0 $X=76560 $Y=339280
X1179 67 11 10 55 87 88 ACHCONX2 $T=108460 188500 0 0 $X=107880 $Y=188140
X1180 821 11 10 796 1619 395 ACHCONX2 $T=137460 230260 1 180 $X=107880 $Y=229900
X1181 802 11 10 806 390 1792 ACHCONX2 $T=108460 261580 0 0 $X=107880 $Y=261220
X1182 1082 11 10 1105 1622 382 ACHCONX2 $T=108460 313780 1 0 $X=107880 $Y=307960
X1183 1081 11 10 1105 1621 393 ACHCONX2 $T=108460 324220 1 0 $X=107880 $Y=318400
X1184 1089 11 10 1097 1625 366 ACHCONX2 $T=108460 334660 1 0 $X=107880 $Y=328840
X1185 821 11 10 797 1620 398 ACHCONX2 $T=109040 219820 0 0 $X=108460 $Y=219460
X1186 812 11 10 1146 418 381 ACHCONX2 $T=109620 282460 1 0 $X=109040 $Y=276640
X1187 803 11 10 806 1626 1791 ACHCONX2 $T=111940 261580 1 0 $X=111360 $Y=255760
X1188 811 11 10 1146 410 1625 ACHCONX2 $T=115420 303340 1 0 $X=114840 $Y=297520
X1189 809 11 10 814 1628 391 ACHCONX2 $T=117160 230260 1 0 $X=116580 $Y=224440
X1190 808 11 10 814 396 1626 ACHCONX2 $T=121800 251140 0 0 $X=121220 $Y=250780
X1191 817 11 10 1109 1777 1421 ACHCONX2 $T=156020 198940 1 180 $X=126440 $Y=198580
X1192 1111 11 10 1142 1723 1627 ACHCONX2 $T=156600 292900 0 180 $X=127020 $Y=287080
X1193 1100 11 10 1177 1405 1725 ACHCONX2 $T=137460 261580 0 0 $X=136880 $Y=261220
X1194 1172 11 10 1112 1407 1727 ACHCONX2 $T=137460 292900 0 0 $X=136880 $Y=292540
X1195 857 11 10 818 1632 396 ACHCONX2 $T=167040 219820 1 180 $X=137460 $Y=219460
X1196 1125 11 10 1118 392 417 ACHCONX2 $T=146160 324220 1 0 $X=145580 $Y=318400
X1197 857 11 10 817 481 1628 ACHCONX2 $T=147320 219820 1 0 $X=146740 $Y=214000
X1198 1125 11 10 1117 382 1629 ACHCONX2 $T=149640 303340 1 0 $X=149060 $Y=297520
X1199 99 11 10 75 109 424 ACHCONX2 $T=154860 188500 0 0 $X=154280 $Y=188140
X1200 1176 11 10 1117 1732 1631 ACHCONX2 $T=161820 272020 1 0 $X=161240 $Y=266200
X1201 1136 11 10 1133 416 434 ACHCONX2 $T=165300 303340 0 0 $X=164720 $Y=302980
X1202 826 11 10 823 398 1630 ACHCONX2 $T=165880 230260 1 0 $X=165300 $Y=224440
X1203 827 11 10 823 394 413 ACHCONX2 $T=194880 240700 1 180 $X=165300 $Y=240340
X1204 820 11 10 1124 1778 1440 ACHCONX2 $T=167040 219820 0 0 $X=166460 $Y=219460
X1205 1162 11 10 1143 479 419 ACHCONX2 $T=167040 282460 1 0 $X=166460 $Y=276640
X1206 1137 11 10 1133 1629 446 ACHCONX2 $T=167040 292900 1 0 $X=166460 $Y=287080
X1207 833 11 10 830 1630 469 ACHCONX2 $T=198360 219820 0 0 $X=197780 $Y=219460
X1208 838 11 10 836 477 476 ACHCONX2 $T=198360 230260 0 0 $X=197780 $Y=229900
X1209 832 11 10 830 412 478 ACHCONX2 $T=198360 240700 0 0 $X=197780 $Y=240340
X1210 1143 11 10 1163 1633 410 ACHCONX2 $T=198360 282460 0 0 $X=197780 $Y=282100
X1211 1169 11 10 1155 445 472 ACHCONX2 $T=198360 292900 0 0 $X=197780 $Y=292540
X1212 835 11 10 838 469 1634 ACHCONX2 $T=200100 240700 1 0 $X=199520 $Y=234880
X1213 1155 11 10 1177 1687 1591 ACHCONX2 $T=229680 261580 0 180 $X=200100 $Y=255760
X1214 1154 11 10 1177 1686 1635 ACHCONX2 $T=204740 272020 1 0 $X=204160 $Y=266200
X1215 1159 11 10 1184 494 480 ACHCONX2 $T=204740 272020 0 0 $X=204160 $Y=271660
X1216 1168 11 10 1155 433 484 ACHCONX2 $T=219240 313780 1 0 $X=218660 $Y=307960
X1217 1123 11 10 847 1737 1632 ACHCONX2 $T=256360 219820 1 180 $X=226780 $Y=219460
X1218 1158 11 10 1184 485 1633 ACHCONX2 $T=227360 282460 0 0 $X=226780 $Y=282100
X1219 848 11 10 871 1636 487 ACHCONX2 $T=235480 240700 1 0 $X=234900 $Y=234880
X1220 847 11 10 871 489 1450 ACHCONX2 $T=237800 261580 1 0 $X=237220 $Y=255760
X1221 1188 11 10 1176 1591 1637 ACHCONX2 $T=238380 272020 1 0 $X=237800 $Y=266200
X1222 859 11 10 862 164 1451 ACHCONX2 $T=239540 219820 1 0 $X=238960 $Y=214000
X1223 1176 11 10 1189 1635 1638 ACHCONX2 $T=240120 282460 1 0 $X=239540 $Y=276640
X1224 1173 11 10 1181 1637 485 ACHCONX2 $T=241280 292900 1 0 $X=240700 $Y=287080
X1225 866 11 10 845 1634 497 ACHCONX2 $T=249980 251140 1 0 $X=249400 $Y=245320
X1226 1173 11 10 1180 1638 495 ACHCONX2 $T=253460 261580 0 0 $X=252880 $Y=261220
X1227 759 11 10 869 496 489 ACHCONX2 $T=283620 251140 1 180 $X=254040 $Y=250780
X1228 153 11 10 162 167 499 ACHCONX2 $T=256940 188500 0 0 $X=256360 $Y=188140
X1229 859 11 10 863 498 500 ACHCONX2 $T=256940 209380 1 0 $X=256360 $Y=203560
X1230 865 11 10 845 475 492 ACHCONX2 $T=256940 219820 0 0 $X=256360 $Y=219460
X1231 759 11 10 868 492 1636 ACHCONX2 $T=256940 230260 1 0 $X=256360 $Y=224440
X1232 1195 11 10 1189 471 1793 ACHCONX2 $T=256940 292900 0 0 $X=256360 $Y=292540
X1233 1194 11 10 1189 483 1794 ACHCONX2 $T=256940 303340 0 0 $X=256360 $Y=302980
X1234 1201 11 10 1180 1794 1639 ACHCONX2 $T=256940 313780 0 0 $X=256360 $Y=313420
X1235 1200 11 10 1180 1793 1640 ACHCONX2 $T=256940 324220 0 0 $X=256360 $Y=323860
X1236 1204 11 10 1185 1640 1553 ACHCONX2 $T=256940 345100 1 0 $X=256360 $Y=339280
X1237 1203 11 10 1185 1639 1552 ACHCONX2 $T=256940 345100 0 0 $X=256360 $Y=344740
X1238 885 11 10 876 526 1453 ACHCONX2 $T=298700 261580 1 0 $X=298120 $Y=255760
X1239 886 11 10 876 1641 520 ACHCONX2 $T=301020 272020 0 0 $X=300440 $Y=271660
X1240 883 11 10 904 1642 526 ACHCONX2 $T=313200 261580 0 0 $X=312620 $Y=261220
X1241 901 11 10 920 1643 541 ACHCONX2 $T=314360 303340 1 0 $X=313780 $Y=297520
X1242 900 11 10 920 1644 531 ACHCONX2 $T=314360 303340 0 0 $X=313780 $Y=302980
X1243 874 11 10 889 557 528 ACHCONX2 $T=314940 230260 0 0 $X=314360 $Y=229900
X1244 897 11 10 175 1739 532 ACHCONX2 $T=317840 198940 0 0 $X=317260 $Y=198580
X1245 959 11 10 913 535 1646 ACHCONX2 $T=317840 345100 1 0 $X=317260 $Y=339280
X1246 903 11 10 883 528 1641 ACHCONX2 $T=348000 251140 1 180 $X=318420 $Y=250780
X1247 888 11 10 874 555 1642 ACHCONX2 $T=319580 230260 1 0 $X=319000 $Y=224440
X1248 910 11 10 1317 1645 533 ACHCONX2 $T=322480 355540 0 0 $X=321900 $Y=355180
X1249 913 11 10 960 533 554 ACHCONX2 $T=323060 334660 0 0 $X=322480 $Y=334300
X1250 909 11 10 1317 1600 536 ACHCONX2 $T=323060 355540 1 0 $X=322480 $Y=349720
X1251 907 11 10 936 1648 1644 ACHCONX2 $T=324220 282460 1 0 $X=323640 $Y=276640
X1252 936 11 10 906 1647 1643 ACHCONX2 $T=324220 282460 0 0 $X=323640 $Y=282100
X1253 210 11 10 206 1779 1458 ACHCONX2 $T=371200 219820 1 180 $X=341620 $Y=219460
X1254 942 11 10 891 541 1462 ACHCONX2 $T=372940 303340 1 180 $X=343360 $Y=302980
X1255 922 11 10 207 1650 558 ACHCONX2 $T=346840 198940 0 0 $X=346260 $Y=198580
X1256 923 11 10 207 1649 555 ACHCONX2 $T=346840 209380 1 0 $X=346260 $Y=203560
X1257 933 11 10 1213 1742 1648 ACHCONX2 $T=346840 272020 0 0 $X=346260 $Y=271660
X1258 891 11 10 943 530 559 ACHCONX2 $T=375840 313780 1 180 $X=346260 $Y=313420
X1259 927 11 10 1209 553 1567 ACHCONX2 $T=346840 334660 1 0 $X=346260 $Y=328840
X1260 928 11 10 1209 1646 1566 ACHCONX2 $T=346840 345100 1 0 $X=346260 $Y=339280
X1261 924 11 10 1286 1740 1645 ACHCONX2 $T=346840 365980 1 0 $X=346260 $Y=360160
X1262 216 11 10 219 1604 1649 ACHCONX2 $T=378160 198940 1 0 $X=377580 $Y=193120
X1263 217 11 10 219 1651 1650 ACHCONX2 $T=378160 198940 0 0 $X=377580 $Y=198580
X1264 1211 11 10 937 1795 573 ACHCONX2 $T=378160 313780 1 0 $X=377580 $Y=307960
X1265 954 11 10 206 1568 1751 ACHCONX2 $T=378740 219820 0 0 $X=378160 $Y=219460
X1266 936 11 10 1211 1781 1477 ACHCONX2 $T=382220 292900 1 0 $X=381640 $Y=287080
X1267 976 11 10 1286 1374 1747 ACHCONX2 $T=382800 365980 1 0 $X=382220 $Y=360160
X1268 229 11 10 227 1488 1748 ACHCONX2 $T=397300 188500 0 0 $X=396720 $Y=188140
X1269 974 11 10 1212 1661 616 ACHCONX2 $T=397880 272020 1 0 $X=397300 $Y=266200
X1270 962 11 10 208 1755 581 ACHCONX2 $T=399620 240700 0 0 $X=399040 $Y=240340
X1271 985 11 10 1317 1756 624 ACHCONX2 $T=400780 334660 0 0 $X=400200 $Y=334300
X1272 959 11 10 1312 1783 1498 ACHCONX2 $T=406000 376420 1 0 $X=405420 $Y=370600
X1273 993 11 10 1212 1757 644 ACHCONX2 $T=418180 240700 1 0 $X=417600 $Y=234880
X1274 991 11 10 219 1759 1652 ACHCONX2 $T=419340 198940 1 0 $X=418760 $Y=193120
X1275 999 11 10 1210 1763 689 ACHCONX2 $T=436740 272020 1 0 $X=436160 $Y=266200
X1276 1014 11 10 1213 1785 1515 ACHCONX2 $T=468060 230260 1 0 $X=467480 $Y=224440
X1277 268 11 10 271 1653 287 ACHCONX2 $T=468060 376420 1 0 $X=467480 $Y=370600
X1278 1023 11 10 1219 1654 1578 ACHCONX2 $T=469220 282460 1 0 $X=468640 $Y=276640
X1279 1035 11 10 1286 1788 1517 ACHCONX2 $T=471540 313780 0 0 $X=470960 $Y=313420
X1280 1024 11 10 1219 1655 1579 ACHCONX2 $T=473860 282460 0 0 $X=473280 $Y=282100
X1281 1026 11 10 1328 1768 1581 ACHCONX2 $T=475020 334660 0 0 $X=474440 $Y=334300
X1282 1213 11 10 261 1796 736 ACHCONX2 $T=475600 219820 0 0 $X=475020 $Y=219460
X1283 276 11 10 274 293 1580 ACHCONX2 $T=479080 198940 1 0 $X=478500 $Y=193120
X1284 1035 11 10 1052 1797 1655 ACHCONX2 $T=492420 292900 0 0 $X=491840 $Y=292540
X1285 1055 11 10 1312 1380 1770 ACHCONX2 $T=495320 345100 0 0 $X=494740 $Y=344740
X1286 1035 11 10 1053 1798 1654 ACHCONX2 $T=499380 282460 1 0 $X=498800 $Y=276640
X1287 1038 11 10 1210 1658 301 ACHCONX2 $T=504020 209380 0 0 $X=503440 $Y=209020
X1288 261 11 10 304 1656 756 ACHCONX2 $T=506920 198940 0 0 $X=506340 $Y=198580
X1289 1040 11 10 1211 1382 1774 ACHCONX2 $T=508080 251140 0 0 $X=507500 $Y=250780
X1290 1039 11 10 1210 1657 1656 ACHCONX2 $T=508660 209380 1 0 $X=508080 $Y=203560
X1291 1066 11 10 1312 1660 1797 ACHCONX2 $T=510400 292900 1 0 $X=509820 $Y=287080
X1292 1065 11 10 1312 1659 1798 ACHCONX2 $T=510980 272020 0 0 $X=510400 $Y=271660
X1293 1062 11 10 1328 1775 1660 ACHCONX2 $T=512140 324220 1 0 $X=511560 $Y=318400
X1294 1346 11 10 561 1349 190 1464 AND4XL $T=365400 240700 1 0 $X=364800 $Y=234880
X1295 574 11 10 588 1469 199 1471 AND4XL $T=389180 303340 0 0 $X=388580 $Y=302980
X1296 1351 11 10 571 592 222 1473 AND4XL $T=393820 355540 1 0 $X=393220 $Y=349720
X1297 1354 11 10 583 602 231 1481 AND4XL $T=404840 261580 0 0 $X=404240 $Y=261220
X1298 1356 11 10 626 1359 198 1487 AND4XL $T=421660 355540 0 180 $X=415840 $Y=349720
X1299 1361 11 10 700 1363 222 1519 AND4XL $T=476760 303340 0 0 $X=476160 $Y=302980
X1300 737 11 10 719 1513 231 1520 AND4XL $T=488940 230260 0 0 $X=488340 $Y=229900
X1301 1364 11 10 748 1522 198 1524 AND4XL $T=505180 334660 1 0 $X=504580 $Y=328840
X1302 1368 11 10 744 741 199 1528 AND4XL $T=509240 251140 1 0 $X=508640 $Y=245320
X1303 27 11 10 767 33 1799 764 ADDFXL $T=48140 365980 1 0 $X=47540 $Y=360160
X1304 1800 11 10 74 71 76 1074 ADDFXL $T=132240 376420 0 180 $X=116560 $Y=370600
X1305 1801 11 10 1122 73 1802 1084 ADDFXL $T=133980 355540 1 180 $X=118300 $Y=355180
X1306 1803 11 10 1116 74 1801 1095 ADDFXL $T=135140 355540 0 180 $X=119460 $Y=349720
X1307 449 11 10 1130 84 1803 1080 ADDFXL $T=145000 345100 1 180 $X=129320 $Y=344740
X1308 1804 11 10 1121 73 1805 1083 ADDFXL $T=145000 365980 0 180 $X=129320 $Y=360160
X1309 1806 11 10 89 85 90 1091 ADDFXL $T=145580 365980 1 180 $X=129900 $Y=365620
X1310 1807 11 10 84 85 1800 1090 ADDFXL $T=147320 376420 0 180 $X=131640 $Y=370600
X1311 1808 11 10 1115 74 1804 1094 ADDFXL $T=149060 355540 1 180 $X=133380 $Y=355180
X1312 420 11 10 1129 84 1808 1079 ADDFXL $T=160080 365980 0 180 $X=144400 $Y=360160
X1313 1805 11 10 1140 100 1809 1127 ADDFXL $T=149060 355540 0 0 $X=148460 $Y=355180
X1314 1802 11 10 1141 100 1810 1128 ADDFXL $T=164140 355540 0 0 $X=163540 $Y=355180
X1315 1810 11 10 1151 68 1811 1139 ADDFXL $T=179220 355540 0 0 $X=178620 $Y=355180
X1316 1809 11 10 1150 68 1812 1138 ADDFXL $T=180960 365980 1 0 $X=180360 $Y=360160
X1317 1813 11 10 1166 121 1806 1149 ADDFXL $T=213440 365980 0 180 $X=197760 $Y=360160
X1318 1814 11 10 1167 121 1807 1148 ADDFXL $T=198940 355540 1 0 $X=198340 $Y=349720
X1319 1815 11 10 1152 1193 1389 1144 ADDFXL $T=230840 324220 1 180 $X=215160 $Y=323860
X1320 1816 11 10 131 142 1814 1164 ADDFXL $T=219240 355540 1 0 $X=218640 $Y=349720
X1321 1817 11 10 134 142 1813 1165 ADDFXL $T=219820 355540 0 0 $X=219220 $Y=355180
X1322 1818 11 10 142 144 1713 1205 ADDFXL $T=229100 365980 0 0 $X=228500 $Y=365620
X1323 1812 11 10 148 120 1819 1170 ADDFXL $T=232580 365980 1 0 $X=231980 $Y=360160
X1324 1820 11 10 1193 146 1816 1186 ADDFXL $T=249400 355540 0 180 $X=233720 $Y=349720
X1325 1811 11 10 152 120 1821 1171 ADDFXL $T=234900 355540 0 0 $X=234300 $Y=355180
X1326 441 11 10 1199 152 1822 1190 ADDFXL $T=237220 334660 0 0 $X=236620 $Y=334300
X1327 1822 11 10 143 157 1820 1182 ADDFXL $T=241860 345100 0 0 $X=241260 $Y=344740
X1328 1823 11 10 146 160 1818 1202 ADDFXL $T=246500 365980 0 0 $X=245900 $Y=365620
X1329 1819 11 10 161 135 151 1196 ADDFXL $T=246500 376420 1 0 $X=245900 $Y=370600
X1330 1821 11 10 157 135 1823 1197 ADDFXL $T=247660 365980 1 0 $X=247060 $Y=360160
X1331 1824 11 10 163 157 1825 1183 ADDFXL $T=264480 355540 0 180 $X=248800 $Y=349720
X1332 1825 11 10 1192 146 1817 1187 ADDFXL $T=265060 355540 1 180 $X=249380 $Y=355180
X1333 435 11 10 1198 152 1824 1191 ADDFXL $T=262740 334660 0 0 $X=262140 $Y=334300
X1334 462 451 11 10 452 61 1826 813 MXI3X1 $T=210540 334660 0 180 $X=197760 $Y=328840
X1335 1317 11 10 1286 29 221 690 691 1782 SDFFRX1 $T=427460 303340 1 0 $X=426860 $Y=297520
X1336 1328 11 10 1312 29 221 690 691 1786 SDFFRX1 $T=444280 292900 0 0 $X=443680 $Y=292540
X1337 1153 91 11 10 1827 1114 XOR3XL $T=137460 313780 1 0 $X=136860 $Y=307960
X1338 91 1121 11 10 1542 1119 XOR3XL $T=165300 345100 1 0 $X=164700 $Y=339280
X1339 114 116 11 10 111 1131 XOR3XL $T=196040 376420 0 180 $X=178040 $Y=370600
X1340 143 1152 11 10 1815 1160 XOR3XL $T=237220 334660 0 180 $X=219220 $Y=328840
X1341 1799 34 11 10 28 NAND2BX1 $T=55680 365980 0 0 $X=55080 $Y=365620
X1342 1537 1828 11 10 1706 NAND2BX1 $T=140360 355540 1 0 $X=139760 $Y=349720
X1343 1789 1431 11 10 1704 NAND2BX1 $T=161820 345100 0 180 $X=157740 $Y=339280
X1344 1596 1193 11 10 1152 NAND2BX1 $T=228520 324220 0 180 $X=224440 $Y=318400
X1345 1790 1596 11 10 1716 NAND2BX1 $T=234320 324220 0 0 $X=233720 $Y=323860
X1346 518 1454 11 10 175 NAND2BX1 $T=317260 209380 1 0 $X=316660 $Y=203560
X1347 1359 1490 11 10 1328 NAND2BX1 $T=423400 355540 0 0 $X=422800 $Y=355180
X1348 1363 1512 11 10 1317 NAND2BX1 $T=479660 303340 1 0 $X=479060 $Y=297520
X1349 39 1532 11 10 1533 1232 MX2X1 $T=97440 345100 1 180 $X=91620 $Y=344740
X1350 37 1791 11 10 1792 1237 MX2X1 $T=114260 251140 0 0 $X=113660 $Y=250780
X1351 39 1794 11 10 1793 1278 MX2X1 $T=275500 292900 1 0 $X=274900 $Y=287080
X1352 39 1552 11 10 1553 1280 MX2X1 $T=277820 334660 0 0 $X=277220 $Y=334300
X1353 198 1566 11 10 1567 1298 MX2X1 $T=365400 334660 0 0 $X=364800 $Y=334300
X1354 199 278 11 10 1580 1332 MX2X1 $T=481980 209380 1 0 $X=481380 $Y=203560
X1355 198 1578 11 10 1579 1330 MX2X1 $T=498220 292900 0 180 $X=492400 $Y=287080
X1356 198 1798 11 10 1797 1343 MX2X1 $T=522000 282460 0 0 $X=521400 $Y=282100
X1357 1584 11 10 1720 794 1109 AOI2BB1X1 $T=96860 219820 1 180 $X=91620 $Y=219460
X1358 1829 11 10 1537 1130 83 AOI2BB1X1 $T=139200 345100 0 180 $X=133960 $Y=339280
X1359 1776 11 10 1828 91 1121 AOI2BB1X1 $T=149640 345100 1 180 $X=144400 $Y=344740
X1360 1665 11 10 1627 1112 408 AOI2BB1X1 $T=146740 282460 0 0 $X=146140 $Y=282100
X1361 1828 11 10 1250 1122 83 AOI2BB1X1 $T=169940 345100 0 0 $X=169340 $Y=344740
X1362 1667 11 10 1631 1177 427 AOI2BB1X1 $T=182120 282460 0 0 $X=181520 $Y=282100
X1363 1668 11 10 1387 827 1124 AOI2BB1X1 $T=184440 209380 0 0 $X=183840 $Y=209020
X1364 1830 11 10 545 1718 1395 AOI2BB1X1 $T=358440 251140 0 0 $X=357840 $Y=250780
X1365 1676 11 10 236 972 206 AOI2BB1X1 $T=417020 209380 1 180 $X=411780 $Y=209020
X1366 666 11 10 1652 227 1571 AOI2BB1X1 $T=450660 209380 0 180 $X=445420 $Y=203560
X1367 675 11 10 1764 1003 1312 AOI2BB1X1 $T=459360 355540 1 0 $X=458760 $Y=349720
X1368 355 11 10 1619 1109 1413 OAI2BB1X1 $T=92220 219820 1 180 $X=87560 $Y=219460
X1369 451 11 10 1390 1442 420 OAI2BB1X1 $T=204160 345100 0 180 $X=199500 $Y=339280
X1370 545 11 10 1394 208 567 OAI2BB1X1 $T=361920 240700 0 0 $X=361320 $Y=240340
X1371 1351 11 10 1601 951 1317 OAI2BB1X1 $T=392080 355540 0 180 $X=387420 $Y=349720
X1372 577 11 10 1647 1212 1467 OAI2BB1X1 $T=394400 272020 0 180 $X=389740 $Y=266200
X1373 1751 11 10 235 971 206 OAI2BB1X1 $T=408320 219820 1 0 $X=407720 $Y=214000
X1374 633 11 10 1383 1211 657 OAI2BB1X1 $T=442540 282460 1 0 $X=441940 $Y=276640
X1375 262 11 10 1611 227 258 OAI2BB1X1 $T=464000 198940 0 180 $X=459340 $Y=193120
X1376 1769 11 10 1659 1312 1526 OAI2BB1X1 $T=508080 324220 1 0 $X=507480 $Y=318400
X1377 1772 11 10 1656 1211 1527 OAI2BB1X1 $T=519100 219820 1 180 $X=514440 $Y=219460
X1378 1831 1703 1627 11 10 NOR2XL $T=103820 282460 0 0 $X=103220 $Y=282100
X1379 1541 1789 1243 11 10 NOR2XL $T=157180 334660 0 180 $X=154260 $Y=328840
X1380 1832 1712 431 11 10 NOR2XL $T=200680 272020 1 180 $X=197760 $Y=271660
X1381 1554 1790 1264 11 10 NOR2XL $T=242440 324220 1 180 $X=239520 $Y=323860
X1382 1830 1692 11 10 INVXL $T=358440 251140 1 180 $X=356100 $Y=250780
X1383 37 11 10 1587 1423 1538 389 NOR4BBX1 $T=133400 209380 0 0 $X=132800 $Y=209020
X1384 54 11 10 1668 1434 1546 454 NOR4BBX1 $T=182120 209380 1 0 $X=181520 $Y=203560
X1385 1427 11 10 1112 1666 AND2X1 $T=151960 282460 1 0 $X=151360 $Y=276640
X1386 1469 11 10 1795 1749 AND2X1 $T=394400 303340 0 0 $X=393800 $Y=302980
X1387 1513 11 10 1796 1766 AND2X1 $T=488940 230260 1 180 $X=484860 $Y=229900
X1388 1087 11 10 69 68 CLKXOR2X1 $T=116000 376420 0 180 $X=109020 $Y=370600
X1389 1826 11 10 1715 1594 CLKXOR2X1 $T=207060 334660 0 0 $X=206460 $Y=334300
X1390 1096 1111 11 10 1722 1831 OAI21X1 $T=101500 292900 0 0 $X=100900 $Y=292540
X1391 1177 1154 11 10 1734 1832 OAI21X1 $T=218080 282460 0 180 $X=214000 $Y=276640
X1392 1559 1271 1598 11 10 1560 NOR3BX1 $T=266800 324220 1 0 $X=266200 $Y=318400
X1393 1829 11 10 1827 1539 1536 NOR3X1 $T=146740 334660 0 0 $X=146140 $Y=334300
.ends MASCO__P2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OAI33XL                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OAI33XL A0 A1 VDD VSS A2 B2 Y B1 B0
** N=14 EP=9 FDC=12
M0 10 A0 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=960 $Y=1080 $dt=0
M1 VSS A1 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1800 $Y=1080 $dt=0
M2 10 A2 VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=2640 $Y=1080 $dt=0
M3 Y B2 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=3480 $Y=1080 $dt=0
M4 10 B1 Y VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=4320 $Y=1080 $dt=0
M5 Y B0 10 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=5160 $Y=1080 $dt=0
M6 11 A0 VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1360 $Y=3600 $dt=1
M7 12 A1 11 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1800 $Y=3600 $dt=1
M8 Y A2 12 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=2640 $Y=3600 $dt=1
M9 13 B2 Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=3480 $Y=3600 $dt=1
M10 14 B1 13 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4320 $Y=3600 $dt=1
M11 VDD B0 14 VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=4760 $Y=3600 $dt=1
.ends OAI33XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2XL                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2XL A Y VDD VSS B
** N=6 EP=5 FDC=4
M0 6 A VSS VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=800 $Y=1360 $dt=0
M1 Y B 6 VSS nmos1v L=1e-07 W=2.4e-07 fw=2.4e-07 simw=2.4e-07 $X=1240 $Y=1360 $dt=0
M2 Y A VDD VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=680 $Y=2760 $dt=1
M3 VDD B Y VDD pmos1v L=1e-07 W=3.6e-07 fw=3.6e-13 simw=3.6e-07 $X=1520 $Y=2760 $dt=1
.ends NAND2XL

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__P3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__P3 2 4 5 7 8 14 15 16 17 18
+ 20 21 22 25 26 27 28 29 30 31
+ 32 33 34 35 36 37 38 39 41 42
+ 43 44 45 46 47 48 49 50 51 52
+ 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72
+ 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92
+ 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112
+ 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132
+ 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152
+ 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172
+ 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192
+ 193 194 195 196 197 198 199 200 201 202
+ 203
** N=1812 EP=191 FDC=23592
X0 204 15 14 21 CLKBUFX2 $T=34800 491260 1 0 $X=34200 $Y=485440
X1 205 15 14 2 CLKBUFX2 $T=36540 459940 0 0 $X=35940 $Y=459580
X2 206 15 14 8 CLKBUFX2 $T=37120 386860 0 0 $X=36520 $Y=386500
X3 207 15 14 7 CLKBUFX2 $T=37120 397300 0 0 $X=36520 $Y=396940
X4 208 15 14 25 CLKBUFX2 $T=37120 512140 0 0 $X=36520 $Y=511780
X5 209 15 14 4 CLKBUFX2 $T=38860 418180 0 0 $X=38260 $Y=417820
X6 210 15 14 22 CLKBUFX2 $T=38860 439060 0 0 $X=38260 $Y=438700
X7 211 15 14 26 CLKBUFX2 $T=40020 543460 0 0 $X=39420 $Y=543100
X8 212 15 14 20 CLKBUFX2 $T=40020 553900 1 0 $X=39420 $Y=548080
X9 213 15 14 29 CLKBUFX2 $T=40600 386860 0 0 $X=40000 $Y=386500
X10 23 15 14 35 CLKBUFX2 $T=51040 376420 0 0 $X=50440 $Y=376060
X11 214 15 14 38 CLKBUFX2 $T=60900 553900 1 0 $X=60300 $Y=548080
X12 215 15 14 17 CLKBUFX2 $T=62060 553900 0 0 $X=61460 $Y=553540
X13 216 15 14 42 CLKBUFX2 $T=81780 553900 1 0 $X=81180 $Y=548080
X14 217 15 14 18 CLKBUFX2 $T=82940 553900 0 0 $X=82340 $Y=553540
X15 218 15 14 52 CLKBUFX2 $T=102660 543460 0 0 $X=102060 $Y=543100
X16 219 15 14 53 CLKBUFX2 $T=102660 553900 1 0 $X=102060 $Y=548080
X17 220 15 14 61 CLKBUFX2 $T=125860 553900 1 0 $X=125260 $Y=548080
X18 221 15 14 60 CLKBUFX2 $T=127020 553900 0 0 $X=126420 $Y=553540
X19 222 15 14 70 CLKBUFX2 $T=147320 553900 1 0 $X=146720 $Y=548080
X20 223 15 14 16 CLKBUFX2 $T=169360 553900 0 0 $X=168760 $Y=553540
X21 224 15 14 55 CLKBUFX2 $T=189660 553900 0 0 $X=189060 $Y=553540
X22 225 15 14 69 CLKBUFX2 $T=191400 553900 1 0 $X=190800 $Y=548080
X23 226 15 14 58 CLKBUFX2 $T=231420 553900 1 0 $X=230820 $Y=548080
X24 227 15 14 100 CLKBUFX2 $T=233160 533020 1 0 $X=232560 $Y=527200
X25 228 15 14 46 CLKBUFX2 $T=251140 553900 0 0 $X=250540 $Y=553540
X26 229 15 14 112 CLKBUFX2 $T=272020 553900 0 0 $X=271420 $Y=553540
X27 230 15 14 113 CLKBUFX2 $T=275500 553900 0 0 $X=274900 $Y=553540
X28 231 15 14 37 CLKBUFX2 $T=288260 553900 1 0 $X=287660 $Y=548080
X29 83 15 14 232 CLKINVX2 $T=198360 407740 0 0 $X=197760 $Y=407380
X30 83 15 14 30 CLKINVX2 $T=201260 407740 0 0 $X=200660 $Y=407380
X31 83 15 14 233 CLKINVX2 $T=213440 397300 0 0 $X=212840 $Y=396940
X32 83 15 14 234 CLKINVX2 $T=397880 418180 0 0 $X=397280 $Y=417820
X33 83 15 14 235 CLKINVX2 $T=400780 418180 0 0 $X=400180 $Y=417820
X34 236 237 15 14 CLKINVX1 $T=179800 397300 1 180 $X=177460 $Y=396940
X35 238 239 15 14 CLKINVX1 $T=185600 386860 0 0 $X=185000 $Y=386500
X36 240 241 15 14 CLKINVX1 $T=213440 470380 0 0 $X=212840 $Y=470020
X37 242 243 15 14 CLKINVX1 $T=217500 459940 1 0 $X=216900 $Y=454120
X38 244 245 15 14 CLKINVX1 $T=254620 470380 0 0 $X=254020 $Y=470020
X39 246 247 15 14 CLKINVX1 $T=255200 480820 1 0 $X=254600 $Y=475000
X40 248 249 15 14 CLKINVX1 $T=277240 407740 1 0 $X=276640 $Y=401920
X41 250 251 15 14 CLKINVX1 $T=289420 397300 1 0 $X=288820 $Y=391480
X42 252 253 15 14 CLKINVX1 $T=330020 470380 0 180 $X=327680 $Y=464560
X43 254 255 15 14 CLKINVX1 $T=332920 522580 0 180 $X=330580 $Y=516760
X44 256 257 15 14 CLKINVX1 $T=337560 512140 1 180 $X=335220 $Y=511780
X45 258 259 15 14 CLKINVX1 $T=338720 470380 1 180 $X=336380 $Y=470020
X46 260 261 15 14 CLKINVX1 $T=341040 480820 1 0 $X=340440 $Y=475000
X47 262 263 15 14 CLKINVX1 $T=344520 407740 0 0 $X=343920 $Y=407380
X48 264 265 15 14 CLKINVX1 $T=346260 522580 0 180 $X=343920 $Y=516760
X49 266 267 15 14 CLKINVX1 $T=346260 522580 1 180 $X=343920 $Y=522220
X50 268 269 15 14 CLKINVX1 $T=346840 397300 1 180 $X=344500 $Y=396940
X51 270 271 15 14 CLKINVX1 $T=350900 407740 0 0 $X=350300 $Y=407380
X52 272 273 15 14 CLKINVX1 $T=353220 397300 1 180 $X=350880 $Y=396940
X53 274 275 15 14 CLKINVX1 $T=352060 491260 1 0 $X=351460 $Y=485440
X54 276 277 15 14 CLKINVX1 $T=357280 418180 0 0 $X=356680 $Y=417820
X55 278 279 15 14 CLKINVX1 $T=367720 533020 0 180 $X=365380 $Y=527200
X56 280 281 15 14 CLKINVX1 $T=366560 459940 1 0 $X=365960 $Y=454120
X57 282 283 15 14 CLKINVX1 $T=368300 480820 1 0 $X=367700 $Y=475000
X58 284 285 15 14 CLKINVX1 $T=371200 543460 1 180 $X=368860 $Y=543100
X59 286 287 15 14 CLKINVX1 $T=371200 553900 0 0 $X=370600 $Y=553540
X60 288 289 15 14 CLKINVX1 $T=372360 418180 1 0 $X=371760 $Y=412360
X61 290 291 15 14 CLKINVX1 $T=373520 459940 1 0 $X=372920 $Y=454120
X62 292 293 15 14 CLKINVX1 $T=378160 470380 0 0 $X=377560 $Y=470020
X63 294 295 15 14 CLKINVX1 $T=383380 407740 0 0 $X=382780 $Y=407380
X64 296 297 15 14 CLKINVX1 $T=385120 407740 1 0 $X=384520 $Y=401920
X65 298 299 15 14 CLKINVX1 $T=388020 470380 0 180 $X=385680 $Y=464560
X66 300 301 15 14 CLKINVX1 $T=391500 470380 1 180 $X=389160 $Y=470020
X67 302 303 15 14 CLKINVX1 $T=392660 480820 1 180 $X=390320 $Y=480460
X68 304 305 15 14 CLKINVX1 $T=394400 428620 0 180 $X=392060 $Y=422800
X69 306 307 15 14 CLKINVX1 $T=396720 501700 0 180 $X=394380 $Y=495880
X70 308 309 15 14 CLKINVX1 $T=399040 407740 0 180 $X=396700 $Y=401920
X71 310 311 15 14 CLKINVX1 $T=397300 533020 1 0 $X=396700 $Y=527200
X72 312 313 15 14 CLKINVX1 $T=397880 501700 1 0 $X=397280 $Y=495880
X73 314 315 15 14 CLKINVX1 $T=400200 459940 0 0 $X=399600 $Y=459580
X74 316 317 15 14 CLKINVX1 $T=404260 491260 0 180 $X=401920 $Y=485440
X75 318 319 15 14 CLKINVX1 $T=404840 501700 1 0 $X=404240 $Y=495880
X76 320 321 15 14 CLKINVX1 $T=404840 533020 1 0 $X=404240 $Y=527200
X77 322 323 15 14 CLKINVX1 $T=406000 480820 1 0 $X=405400 $Y=475000
X78 324 325 15 14 CLKINVX1 $T=408900 459940 1 0 $X=408300 $Y=454120
X79 326 327 15 14 CLKINVX1 $T=408900 522580 0 0 $X=408300 $Y=522220
X80 328 329 15 14 CLKINVX1 $T=412380 449500 0 180 $X=410040 $Y=443680
X81 330 331 15 14 CLKINVX1 $T=413540 553900 0 180 $X=411200 $Y=548080
X82 332 333 15 14 CLKINVX1 $T=412960 407740 0 0 $X=412360 $Y=407380
X83 334 335 15 14 CLKINVX1 $T=414700 418180 0 180 $X=412360 $Y=412360
X84 336 337 15 14 CLKINVX1 $T=412960 428620 0 0 $X=412360 $Y=428260
X85 338 339 15 14 CLKINVX1 $T=417020 428620 1 180 $X=414680 $Y=428260
X86 340 341 15 14 CLKINVX1 $T=417020 543460 0 180 $X=414680 $Y=537640
X87 342 343 15 14 CLKINVX1 $T=418180 491260 1 180 $X=415840 $Y=490900
X88 344 345 15 14 CLKINVX1 $T=417020 397300 0 0 $X=416420 $Y=396940
X89 346 347 15 14 CLKINVX1 $T=424560 480820 0 0 $X=423960 $Y=480460
X90 348 349 15 14 CLKINVX1 $T=430360 543460 1 180 $X=428020 $Y=543100
X91 350 351 15 14 CLKINVX1 $T=433260 501700 0 180 $X=430920 $Y=495880
X92 352 353 15 14 CLKINVX1 $T=433260 397300 1 0 $X=432660 $Y=391480
X93 354 355 15 14 CLKINVX1 $T=433260 418180 0 0 $X=432660 $Y=417820
X94 356 357 15 14 CLKINVX1 $T=437320 522580 1 180 $X=434980 $Y=522220
X95 358 359 15 14 CLKINVX1 $T=439060 470380 1 180 $X=436720 $Y=470020
X96 360 361 15 14 CLKINVX1 $T=440800 522580 0 0 $X=440200 $Y=522220
X97 362 363 15 14 CLKINVX1 $T=443700 428620 1 0 $X=443100 $Y=422800
X98 364 365 15 14 CLKINVX1 $T=446020 439060 1 180 $X=443680 $Y=438700
X99 366 367 15 14 CLKINVX1 $T=448340 491260 0 180 $X=446000 $Y=485440
X100 368 369 15 14 CLKINVX1 $T=450080 480820 0 180 $X=447740 $Y=475000
X101 370 371 15 14 CLKINVX1 $T=450660 491260 0 180 $X=448320 $Y=485440
X102 372 373 15 14 CLKINVX1 $T=451820 501700 1 180 $X=449480 $Y=501340
X103 374 375 15 14 CLKINVX1 $T=452980 418180 0 180 $X=450640 $Y=412360
X104 376 377 15 14 CLKINVX1 $T=452980 439060 1 180 $X=450640 $Y=438700
X105 378 379 15 14 CLKINVX1 $T=454140 418180 1 180 $X=451800 $Y=417820
X106 380 381 15 14 CLKINVX1 $T=455300 501700 1 180 $X=452960 $Y=501340
X107 382 383 15 14 CLKINVX1 $T=457040 428620 0 180 $X=454700 $Y=422800
X108 384 385 15 14 CLKINVX1 $T=457040 439060 1 180 $X=454700 $Y=438700
X109 386 387 15 14 CLKINVX1 $T=459940 543460 0 180 $X=457600 $Y=537640
X110 388 389 15 14 CLKINVX1 $T=462840 501700 1 180 $X=460500 $Y=501340
X111 390 391 15 14 CLKINVX1 $T=465740 480820 0 180 $X=463400 $Y=475000
X112 392 393 15 14 CLKINVX1 $T=469800 522580 1 180 $X=467460 $Y=522220
X113 394 395 15 14 CLKINVX1 $T=469220 407740 1 0 $X=468620 $Y=401920
X114 396 397 15 14 CLKINVX1 $T=474440 459940 1 0 $X=473840 $Y=454120
X115 398 399 15 14 CLKINVX1 $T=477920 386860 1 0 $X=477320 $Y=381040
X116 400 401 15 14 CLKINVX1 $T=492420 439060 1 180 $X=490080 $Y=438700
X117 402 403 15 14 CLKINVX1 $T=492420 480820 1 0 $X=491820 $Y=475000
X118 404 405 15 14 CLKINVX1 $T=493580 407740 0 0 $X=492980 $Y=407380
X119 406 181 15 14 CLKINVX1 $T=498800 376420 1 180 $X=496460 $Y=376060
X120 407 408 15 14 CLKINVX1 $T=501700 480820 1 180 $X=499360 $Y=480460
X121 409 410 15 14 CLKINVX1 $T=502280 522580 1 180 $X=499940 $Y=522220
X122 411 412 15 14 CLKINVX1 $T=505180 522580 0 180 $X=502840 $Y=516760
X123 413 414 15 14 CLKINVX1 $T=505760 386860 1 0 $X=505160 $Y=381040
X124 415 416 15 14 CLKINVX1 $T=506340 470380 1 0 $X=505740 $Y=464560
X125 417 418 15 14 CLKINVX1 $T=508660 386860 0 0 $X=508060 $Y=386500
X126 419 420 15 14 CLKINVX1 $T=510980 480820 0 180 $X=508640 $Y=475000
X127 421 422 15 14 CLKINVX1 $T=511560 533020 0 180 $X=509220 $Y=527200
X128 423 424 15 14 CLKINVX1 $T=510400 449500 1 0 $X=509800 $Y=443680
X129 425 426 15 14 CLKINVX1 $T=513300 407740 1 180 $X=510960 $Y=407380
X130 427 428 15 14 CLKINVX1 $T=514460 449500 0 0 $X=513860 $Y=449140
X131 429 430 15 14 CLKINVX1 $T=515620 397300 0 0 $X=515020 $Y=396940
X132 431 432 15 14 CLKINVX1 $T=519100 491260 0 180 $X=516760 $Y=485440
X133 433 434 15 14 CLKINVX1 $T=519680 407740 1 180 $X=517340 $Y=407380
X134 435 436 15 14 CLKINVX1 $T=519680 407740 0 0 $X=519080 $Y=407380
X135 437 5 15 14 30 23 DFFRHQX1 $T=51040 376420 1 180 $X=34780 $Y=376060
X136 34 5 15 14 30 207 DFFRHQX1 $T=51040 386860 0 180 $X=34780 $Y=381040
X137 122 5 15 14 233 438 DFFRHQX1 $T=316100 553900 0 180 $X=299840 $Y=548080
X138 123 5 15 14 233 439 DFFRHQX1 $T=316680 553900 1 180 $X=300420 $Y=553540
X139 119 5 15 14 233 440 DFFRHQX1 $T=301600 543460 1 0 $X=301000 $Y=537640
X140 120 5 15 14 233 441 DFFRHQX1 $T=316100 543460 0 0 $X=315500 $Y=543100
X141 124 5 15 14 233 442 DFFRHQX1 $T=319580 553900 1 0 $X=318980 $Y=548080
X142 130 5 15 14 233 443 DFFRHQX1 $T=335820 553900 1 180 $X=319560 $Y=553540
X143 128 5 15 14 233 444 DFFRHQX1 $T=336400 553900 0 0 $X=335800 $Y=553540
X144 132 5 15 14 233 445 DFFRHQX1 $T=337560 553900 1 0 $X=336960 $Y=548080
X145 144 5 15 14 235 446 DFFRHQX1 $T=378160 553900 1 0 $X=377560 $Y=548080
X146 145 5 15 14 235 447 DFFRHQX1 $T=378740 543460 0 0 $X=378140 $Y=543100
X147 146 5 15 14 235 448 DFFRHQX1 $T=383960 553900 0 0 $X=383360 $Y=553540
X148 148 5 15 14 235 449 DFFRHQX1 $T=393820 553900 1 0 $X=393220 $Y=548080
X149 142 5 15 14 235 450 DFFRHQX1 $T=418760 553900 0 0 $X=418160 $Y=553540
X150 152 5 15 14 235 451 DFFRHQX1 $T=434420 553900 1 0 $X=433820 $Y=548080
X151 147 5 15 14 235 452 DFFRHQX1 $T=434420 553900 0 0 $X=433820 $Y=553540
X152 173 5 15 14 235 453 DFFRHQX1 $T=465740 553900 0 180 $X=449480 $Y=548080
X153 174 5 15 14 235 454 DFFRHQX1 $T=465740 553900 1 180 $X=449480 $Y=553540
X154 455 5 15 14 235 456 DFFRHQX1 $T=468060 501700 0 0 $X=467460 $Y=501340
X155 143 5 15 14 235 457 DFFRHQX1 $T=472120 553900 1 0 $X=471520 $Y=548080
X156 458 5 15 14 234 459 DFFRHQX1 $T=473280 439060 0 0 $X=472680 $Y=438700
X157 154 5 15 14 235 460 DFFRHQX1 $T=488940 553900 1 180 $X=472680 $Y=553540
X158 461 5 15 14 235 462 DFFRHQX1 $T=486040 501700 0 0 $X=485440 $Y=501340
X159 177 5 15 14 235 463 DFFRHQX1 $T=488940 553900 1 0 $X=488340 $Y=548080
X160 180 5 15 14 235 464 DFFRHQX1 $T=490100 553900 0 0 $X=489500 $Y=553540
X161 188 5 15 14 235 465 DFFRHQX1 $T=506920 553900 1 0 $X=506320 $Y=548080
X162 184 5 15 14 235 466 DFFRHQX1 $T=506920 553900 0 0 $X=506320 $Y=553540
X163 200 5 15 14 235 467 DFFRHQX1 $T=523740 553900 0 0 $X=523140 $Y=553540
X164 201 5 15 14 235 468 DFFRHQX1 $T=524320 553900 1 0 $X=523720 $Y=548080
X165 469 5 15 14 30 470 471 27 SDFFRHQX1 $T=80620 418180 0 180 $X=60880 $Y=412360
X166 472 5 15 14 30 473 474 27 SDFFRHQX1 $T=81200 397300 1 180 $X=61460 $Y=396940
X167 475 5 15 14 30 476 477 27 SDFFRHQX1 $T=81200 407740 0 180 $X=61460 $Y=401920
X168 478 5 15 14 232 479 480 39 SDFFRHQX1 $T=81780 480820 0 180 $X=62040 $Y=475000
X169 481 5 15 14 232 482 483 39 SDFFRHQX1 $T=63220 459940 1 0 $X=62620 $Y=454120
X170 484 5 15 14 232 485 486 39 SDFFRHQX1 $T=82360 491260 1 180 $X=62620 $Y=490900
X171 487 5 15 14 30 488 489 39 SDFFRHQX1 $T=82940 449500 1 180 $X=63200 $Y=449140
X172 490 5 15 14 30 491 491 27 SDFFRHQX1 $T=83520 386860 1 180 $X=63780 $Y=386500
X173 492 5 15 14 30 493 493 27 SDFFRHQX1 $T=66700 386860 1 0 $X=66100 $Y=381040
X174 494 5 15 14 30 495 495 39 SDFFRHQX1 $T=91060 439060 1 180 $X=71320 $Y=438700
X175 496 5 15 14 232 497 498 39 SDFFRHQX1 $T=96860 439060 0 180 $X=77120 $Y=433240
X176 499 5 15 14 232 500 501 39 SDFFRHQX1 $T=100920 470380 1 180 $X=81180 $Y=470020
X177 502 5 15 14 30 503 504 43 SDFFRHQX1 $T=103820 428620 1 180 $X=84080 $Y=428260
X178 54 5 15 14 30 505 505 45 SDFFRHQX1 $T=105560 386860 1 180 $X=85820 $Y=386500
X179 506 5 15 14 30 507 508 45 SDFFRHQX1 $T=86420 397300 0 0 $X=85820 $Y=396940
X180 509 5 15 14 30 510 510 39 SDFFRHQX1 $T=105560 418180 1 180 $X=85820 $Y=417820
X181 511 5 15 14 30 512 513 43 SDFFRHQX1 $T=105560 428620 0 180 $X=85820 $Y=422800
X182 514 5 15 14 30 515 515 43 SDFFRHQX1 $T=106140 407740 0 180 $X=86400 $Y=401920
X183 516 5 15 14 232 517 518 43 SDFFRHQX1 $T=108460 459940 1 0 $X=107860 $Y=454120
X184 519 5 15 14 30 520 521 45 SDFFRHQX1 $T=129920 407740 0 180 $X=110180 $Y=401920
X185 522 5 15 14 30 523 524 43 SDFFRHQX1 $T=129920 439060 0 180 $X=110180 $Y=433240
X186 525 5 15 14 30 526 527 43 SDFFRHQX1 $T=132820 439060 1 180 $X=113080 $Y=438700
X187 59 5 15 14 30 528 529 45 SDFFRHQX1 $T=134560 397300 1 180 $X=114820 $Y=396940
X188 530 5 15 14 30 531 532 43 SDFFRHQX1 $T=116000 449500 0 0 $X=115400 $Y=449140
X189 533 5 15 14 30 534 535 43 SDFFRHQX1 $T=123540 449500 1 0 $X=122940 $Y=443680
X190 64 5 15 14 30 536 537 45 SDFFRHQX1 $T=149060 407740 0 180 $X=129320 $Y=401920
X191 538 5 15 14 30 539 539 43 SDFFRHQX1 $T=150800 439060 0 180 $X=131060 $Y=433240
X192 540 5 15 14 232 541 542 43 SDFFRHQX1 $T=135140 449500 0 0 $X=134540 $Y=449140
X193 56 5 15 14 30 543 544 45 SDFFRHQX1 $T=157760 407740 0 0 $X=157160 $Y=407380
X194 71 5 15 14 30 545 546 45 SDFFRHQX1 $T=157760 418180 1 0 $X=157160 $Y=412360
X195 77 5 15 14 30 547 548 45 SDFFRHQX1 $T=176900 407740 0 0 $X=176300 $Y=407380
X196 89 5 15 14 30 549 550 45 SDFFRHQX1 $T=217500 418180 1 180 $X=197760 $Y=417820
X197 91 5 15 14 30 551 552 45 SDFFRHQX1 $T=217500 428620 0 180 $X=197760 $Y=422800
X198 134 5 15 14 233 553 554 555 SDFFRHQX1 $T=339880 533020 0 0 $X=339280 $Y=532660
X199 137 5 15 14 233 287 286 556 SDFFRHQX1 $T=352060 553900 0 0 $X=351460 $Y=553540
X200 138 5 15 14 233 285 284 557 SDFFRHQX1 $T=355540 553900 1 0 $X=354940 $Y=548080
X201 121 5 15 14 235 330 331 341 SDFFRHQX1 $T=399620 553900 0 0 $X=399020 $Y=553540
X202 153 5 15 14 235 340 341 558 SDFFRHQX1 $T=401360 543460 0 0 $X=400760 $Y=543100
X203 118 5 15 14 235 349 348 559 SDFFRHQX1 $T=415280 553900 1 0 $X=414680 $Y=548080
X204 560 5 15 14 234 376 377 561 SDFFRHQX1 $T=438480 459940 1 0 $X=437880 $Y=454120
X205 168 5 15 14 235 562 563 564 SDFFRHQX1 $T=446600 522580 1 0 $X=446000 $Y=516760
X206 565 15 14 566 5 30 206 DFFRX1 $T=52200 397300 0 180 $X=34780 $Y=391480
X207 567 15 14 568 5 232 204 DFFRX1 $T=55100 491260 0 180 $X=37680 $Y=485440
X208 569 15 14 570 5 232 205 DFFRX1 $T=56840 459940 1 180 $X=39420 $Y=459580
X209 571 15 14 572 5 232 208 DFFRX1 $T=57420 512140 1 180 $X=40000 $Y=511780
X210 573 15 14 574 5 30 209 DFFRX1 $T=59160 418180 1 180 $X=41740 $Y=417820
X211 575 15 14 576 5 30 213 DFFRX1 $T=59160 439060 0 180 $X=41740 $Y=433240
X212 577 15 14 578 5 30 210 DFFRX1 $T=59160 439060 1 180 $X=41740 $Y=438700
X213 579 15 14 580 5 232 211 DFFRX1 $T=60320 543460 1 180 $X=42900 $Y=543100
X214 581 15 14 582 5 232 212 DFFRX1 $T=60320 553900 0 180 $X=42900 $Y=548080
X215 583 15 14 584 5 232 214 DFFRX1 $T=81200 553900 0 180 $X=63780 $Y=548080
X216 585 15 14 586 5 232 215 DFFRX1 $T=82360 553900 1 180 $X=64940 $Y=553540
X217 587 15 14 588 5 232 216 DFFRX1 $T=102080 553900 0 180 $X=84660 $Y=548080
X218 589 15 14 590 5 232 217 DFFRX1 $T=103240 553900 1 180 $X=85820 $Y=553540
X219 591 15 14 592 5 232 219 DFFRX1 $T=125860 553900 0 180 $X=108440 $Y=548080
X220 593 15 14 594 5 232 218 DFFRX1 $T=127020 553900 1 180 $X=109600 $Y=553540
X221 595 15 14 596 5 232 220 DFFRX1 $T=146160 553900 0 180 $X=128740 $Y=548080
X222 597 15 14 598 5 232 221 DFFRX1 $T=147320 553900 1 180 $X=129900 $Y=553540
X223 599 15 14 600 5 232 222 DFFRX1 $T=167620 553900 0 180 $X=150200 $Y=548080
X224 601 15 14 602 5 232 223 DFFRX1 $T=152540 553900 0 0 $X=151940 $Y=553540
X225 603 15 14 604 5 233 224 DFFRX1 $T=172840 553900 0 0 $X=172240 $Y=553540
X226 605 15 14 606 5 233 225 DFFRX1 $T=174580 553900 1 0 $X=173980 $Y=548080
X227 607 15 14 608 5 233 227 DFFRX1 $T=198360 553900 0 0 $X=197760 $Y=553540
X228 609 15 14 610 5 233 226 DFFRX1 $T=215180 553900 0 0 $X=214580 $Y=553540
X229 611 15 14 612 5 233 228 DFFRX1 $T=234320 553900 0 0 $X=233720 $Y=553540
X230 613 15 14 614 5 233 229 DFFRX1 $T=252300 553900 1 0 $X=251700 $Y=548080
X231 615 15 14 616 5 233 230 DFFRX1 $T=255200 553900 0 0 $X=254600 $Y=553540
X232 617 15 14 618 5 233 231 DFFRX1 $T=269120 553900 1 0 $X=268520 $Y=548080
X233 619 15 14 620 5 233 621 DFFRX1 $T=300440 501700 1 0 $X=299840 $Y=495880
X234 622 15 14 623 5 233 624 DFFRX1 $T=317840 501700 1 180 $X=300420 $Y=501340
X235 625 15 14 626 5 233 627 DFFRX1 $T=327700 449500 1 180 $X=310280 $Y=449140
X236 628 15 14 629 5 233 630 DFFRX1 $T=311460 449500 1 0 $X=310860 $Y=443680
X237 631 15 14 632 5 97 127 DFFRX1 $T=313200 386860 1 0 $X=312600 $Y=381040
X238 633 15 14 634 5 97 131 DFFRX1 $T=317840 376420 0 0 $X=317240 $Y=376060
X239 635 15 14 636 5 233 637 DFFRX1 $T=319580 501700 1 0 $X=318980 $Y=495880
X240 638 15 14 639 5 234 640 DFFRX1 $T=320160 439060 1 0 $X=319560 $Y=433240
X241 641 15 14 642 5 233 643 DFFRX1 $T=320160 501700 0 0 $X=319560 $Y=501340
X242 644 15 14 645 5 97 136 DFFRX1 $T=330020 386860 1 0 $X=329420 $Y=381040
X243 646 15 14 647 5 234 133 DFFRX1 $T=353220 376420 1 180 $X=335800 $Y=376060
X244 648 15 14 649 5 233 650 DFFRX1 $T=338140 501700 0 0 $X=337540 $Y=501340
X245 651 15 14 652 5 233 653 DFFRX1 $T=338720 533020 1 0 $X=338120 $Y=527200
X246 654 15 14 655 5 234 656 DFFRX1 $T=341040 439060 1 0 $X=340440 $Y=433240
X247 657 15 14 658 5 234 659 DFFRX1 $T=341040 470380 1 0 $X=340440 $Y=464560
X248 660 15 14 661 5 234 662 DFFRX1 $T=344520 470380 0 0 $X=343920 $Y=470020
X249 663 15 14 664 5 234 665 DFFRX1 $T=354380 439060 0 0 $X=353780 $Y=438700
X250 666 15 14 667 5 234 668 DFFRX1 $T=354380 512140 0 0 $X=353780 $Y=511780
X251 554 15 14 553 5 234 669 DFFRX1 $T=355540 501700 0 0 $X=354940 $Y=501340
X252 670 15 14 671 5 234 672 DFFRX1 $T=356700 512140 1 0 $X=356100 $Y=506320
X253 673 15 14 674 5 234 140 DFFRX1 $T=357860 376420 0 0 $X=357260 $Y=376060
X254 675 15 14 676 5 234 141 DFFRX1 $T=359020 397300 0 0 $X=358420 $Y=396940
X255 677 15 14 678 5 234 139 DFFRX1 $T=359020 407740 1 0 $X=358420 $Y=401920
X256 679 15 14 680 5 234 681 DFFRX1 $T=375840 522580 0 180 $X=358420 $Y=516760
X257 682 15 14 683 5 234 684 DFFRX1 $T=378160 439060 0 0 $X=377560 $Y=438700
X258 685 15 14 686 5 234 687 DFFRX1 $T=378160 459940 0 0 $X=377560 $Y=459580
X259 688 15 14 689 5 234 690 DFFRX1 $T=378160 512140 0 0 $X=377560 $Y=511780
X260 691 15 14 692 5 234 149 DFFRX1 $T=380480 376420 0 0 $X=379880 $Y=376060
X261 693 15 14 694 5 234 151 DFFRX1 $T=380480 397300 0 0 $X=379880 $Y=396940
X262 695 15 14 696 5 234 697 DFFRX1 $T=380480 512140 1 0 $X=379880 $Y=506320
X263 698 15 14 699 5 234 150 DFFRX1 $T=381060 397300 1 0 $X=380460 $Y=391480
X264 700 15 14 701 5 234 702 DFFRX1 $T=381640 459940 1 0 $X=381040 $Y=454120
X265 703 15 14 704 5 234 705 DFFRX1 $T=387440 449500 0 0 $X=386840 $Y=449140
X266 706 15 14 707 5 234 708 DFFRX1 $T=388020 449500 1 0 $X=387420 $Y=443680
X267 709 15 14 710 5 234 155 DFFRX1 $T=393820 386860 0 0 $X=393220 $Y=386500
X268 711 15 14 712 5 235 713 DFFRX1 $T=411800 512140 1 180 $X=394380 $Y=511780
X269 714 15 14 555 5 235 715 DFFRX1 $T=401360 512140 1 0 $X=400760 $Y=506320
X270 716 15 14 717 5 234 156 DFFRX1 $T=401940 386860 1 0 $X=401340 $Y=381040
X271 718 15 14 719 5 234 157 DFFRX1 $T=404260 376420 0 0 $X=403660 $Y=376060
X272 720 15 14 721 5 234 159 DFFRX1 $T=410640 386860 0 0 $X=410040 $Y=386500
X273 722 15 14 723 5 234 724 DFFRX1 $T=414120 449500 1 0 $X=413520 $Y=443680
X274 725 15 14 726 5 235 727 DFFRX1 $T=419340 522580 1 0 $X=418740 $Y=516760
X275 728 15 14 564 5 235 729 DFFRX1 $T=437320 512140 0 180 $X=419900 $Y=506320
X276 730 15 14 731 5 234 732 DFFRX1 $T=421660 459940 1 0 $X=421060 $Y=454120
X277 733 15 14 734 5 234 735 DFFRX1 $T=422820 459940 0 0 $X=422220 $Y=459580
X278 736 15 14 737 5 234 163 DFFRX1 $T=427460 386860 0 0 $X=426860 $Y=386500
X279 738 15 14 739 5 235 740 DFFRX1 $T=448920 512140 1 180 $X=431500 $Y=511780
X280 741 15 14 742 5 234 167 DFFRX1 $T=454720 397300 0 180 $X=437300 $Y=391480
X281 743 15 14 744 5 234 745 DFFRX1 $T=439640 459940 0 0 $X=439040 $Y=459580
X282 746 15 14 747 5 234 748 DFFRX1 $T=463420 449500 1 180 $X=446000 $Y=449140
X283 749 15 14 750 5 235 751 DFFRX1 $T=447760 470380 1 0 $X=447160 $Y=464560
X284 752 15 14 753 5 165 170 DFFRX1 $T=448920 386860 1 0 $X=448320 $Y=381040
X285 754 15 14 755 5 234 171 DFFRX1 $T=448920 386860 0 0 $X=448320 $Y=386500
X286 756 15 14 757 5 234 172 DFFRX1 $T=448920 397300 0 0 $X=448320 $Y=396940
X287 563 15 14 562 5 235 758 DFFRX1 $T=465740 512140 1 180 $X=448320 $Y=511780
X288 759 15 14 760 5 234 178 DFFRX1 $T=468060 397300 0 0 $X=467460 $Y=396940
X289 761 15 14 762 5 235 763 DFFRX1 $T=468060 470380 1 0 $X=467460 $Y=464560
X290 764 15 14 765 5 235 766 DFFRX1 $T=468640 512140 1 0 $X=468040 $Y=506320
X291 767 15 14 768 5 235 769 DFFRX1 $T=472700 512140 0 0 $X=472100 $Y=511780
X292 770 15 14 771 5 235 772 DFFRX1 $T=476180 459940 1 0 $X=475580 $Y=454120
X293 773 15 14 774 5 234 775 DFFRX1 $T=498800 439060 0 180 $X=481380 $Y=433240
X294 776 15 14 777 5 234 182 DFFRX1 $T=484880 397300 0 0 $X=484280 $Y=396940
X295 778 15 14 779 5 235 780 DFFRX1 $T=484880 470380 1 0 $X=484280 $Y=464560
X296 781 15 14 782 5 165 185 DFFRX1 $T=485460 386860 0 0 $X=484860 $Y=386500
X297 783 15 14 784 5 235 785 DFFRX1 $T=487780 512140 1 0 $X=487180 $Y=506320
X298 786 15 14 787 5 235 788 DFFRX1 $T=490680 512140 0 0 $X=490080 $Y=511780
X299 789 15 14 790 5 165 190 DFFRX1 $T=493000 397300 1 0 $X=492400 $Y=391480
X300 791 15 14 792 5 235 793 DFFRX1 $T=493000 459940 1 0 $X=492400 $Y=454120
X301 794 15 14 795 5 235 796 DFFRX1 $T=505180 501700 0 0 $X=504580 $Y=501340
X302 797 15 14 798 5 235 195 DFFRX1 $T=505180 512140 1 0 $X=504580 $Y=506320
X303 799 15 14 800 5 235 801 DFFRX1 $T=509820 459940 1 0 $X=509220 $Y=454120
X304 802 15 14 803 5 235 804 DFFRX1 $T=522000 449500 0 0 $X=521400 $Y=449140
X305 805 15 14 806 5 235 807 DFFRX1 $T=522000 512140 1 0 $X=521400 $Y=506320
X306 808 15 14 809 5 235 810 DFFRX1 $T=522580 512140 0 0 $X=521980 $Y=511780
X307 811 15 14 812 5 235 813 DFFRX1 $T=523160 522580 1 0 $X=522560 $Y=516760
X308 814 15 14 815 5 235 816 DFFRX1 $T=526640 459940 1 0 $X=526040 $Y=454120
X309 817 15 14 818 5 235 819 DFFRX1 $T=528960 470380 1 0 $X=528360 $Y=464560
X310 820 15 14 821 5 30 822 27 823 SDFFRXL $T=61480 449500 0 180 $X=40000 $Y=443680
X311 824 15 14 825 5 232 826 27 827 SDFFRXL $T=61480 470380 0 180 $X=40000 $Y=464560
X312 828 15 14 829 5 232 830 27 831 SDFFRXL $T=61480 491260 1 180 $X=40000 $Y=490900
X313 832 15 14 833 5 232 834 27 835 SDFFRXL $T=63220 512140 0 180 $X=41740 $Y=506320
X314 836 15 14 837 5 232 838 27 839 SDFFRXL $T=73660 522580 0 180 $X=52180 $Y=516760
X315 840 15 14 841 5 30 842 27 843 SDFFRXL $T=81780 428620 0 180 $X=60300 $Y=422800
X316 844 15 14 845 5 232 846 27 847 SDFFRXL $T=63800 512140 0 0 $X=63200 $Y=511780
X317 848 15 14 849 5 232 850 27 851 SDFFRXL $T=63800 522580 0 0 $X=63200 $Y=522220
X318 852 15 14 853 5 232 854 39 855 SDFFRXL $T=102660 480820 0 180 $X=81180 $Y=475000
X319 44 15 14 856 5 30 857 51 858 SDFFRXL $T=83520 376420 0 0 $X=82920 $Y=376060
X320 859 15 14 860 5 232 861 39 862 SDFFRXL $T=106140 480820 1 180 $X=84660 $Y=480460
X321 863 15 14 864 5 232 865 39 866 SDFFRXL $T=106140 491260 0 180 $X=84660 $Y=485440
X322 867 15 14 868 5 232 869 39 870 SDFFRXL $T=85260 491260 0 0 $X=84660 $Y=490900
X323 871 15 14 872 5 232 873 27 874 SDFFRXL $T=85260 522580 1 0 $X=84660 $Y=516760
X324 875 15 14 876 5 232 877 27 878 SDFFRXL $T=85260 522580 0 0 $X=84660 $Y=522220
X325 879 15 14 880 5 232 881 27 882 SDFFRXL $T=108460 522580 0 0 $X=107860 $Y=522220
X326 883 15 14 884 5 232 885 27 886 SDFFRXL $T=129920 522580 0 180 $X=108440 $Y=516760
X327 887 15 14 888 5 232 889 39 890 SDFFRXL $T=109620 491260 0 0 $X=109020 $Y=490900
X328 891 15 14 892 5 30 893 43 894 SDFFRXL $T=110780 428620 0 0 $X=110180 $Y=428260
X329 895 15 14 896 5 232 897 39 898 SDFFRXL $T=114260 491260 1 0 $X=113660 $Y=485440
X330 899 15 14 900 5 232 901 27 902 SDFFRXL $T=149640 533020 0 180 $X=128160 $Y=527200
X331 903 15 14 904 5 232 905 27 906 SDFFRXL $T=129340 522580 0 0 $X=128740 $Y=522220
X332 907 15 14 908 5 232 909 39 910 SDFFRXL $T=131080 480820 0 0 $X=130480 $Y=480460
X333 911 15 14 912 5 30 913 43 914 SDFFRXL $T=131660 428620 1 0 $X=131060 $Y=422800
X334 915 15 14 916 5 232 917 39 918 SDFFRXL $T=133400 491260 0 0 $X=132800 $Y=490900
X335 919 15 14 920 5 232 921 39 922 SDFFRXL $T=135140 491260 1 0 $X=134540 $Y=485440
X336 923 15 14 924 5 30 925 43 926 SDFFRXL $T=136300 439060 0 0 $X=135700 $Y=438700
X337 927 15 14 48 5 30 928 45 929 SDFFRXL $T=136880 397300 0 0 $X=136280 $Y=396940
X338 930 15 14 57 5 30 931 45 932 SDFFRXL $T=137460 386860 0 0 $X=136860 $Y=386500
X339 67 15 14 68 5 30 933 45 934 SDFFRXL $T=138620 376420 0 0 $X=138020 $Y=376060
X340 935 15 14 65 5 30 936 45 937 SDFFRXL $T=138620 386860 1 0 $X=138020 $Y=381040
X341 938 15 14 939 5 232 940 27 941 SDFFRXL $T=149640 533020 1 0 $X=149040 $Y=527200
X342 942 15 14 943 5 232 944 27 945 SDFFRXL $T=150220 522580 0 0 $X=149620 $Y=522220
X343 946 15 14 947 5 30 948 43 949 SDFFRXL $T=150800 449500 1 0 $X=150200 $Y=443680
X344 950 15 14 951 5 30 952 43 953 SDFFRXL $T=154280 449500 0 0 $X=153680 $Y=449140
X345 954 15 14 955 5 232 956 39 957 SDFFRXL $T=154280 491260 0 0 $X=153680 $Y=490900
X346 958 15 14 959 5 232 960 39 961 SDFFRXL $T=156020 491260 1 0 $X=155420 $Y=485440
X347 962 15 14 963 5 233 964 39 965 SDFFRXL $T=191980 501700 0 180 $X=170500 $Y=495880
X348 966 15 14 967 5 233 968 27 969 SDFFRXL $T=171100 522580 0 0 $X=170500 $Y=522220
X349 970 15 14 971 5 233 972 27 973 SDFFRXL $T=171100 533020 1 0 $X=170500 $Y=527200
X350 974 15 14 975 5 233 976 39 977 SDFFRXL $T=172840 480820 0 0 $X=172240 $Y=480460
X351 978 15 14 979 5 233 980 43 981 SDFFRXL $T=194300 459940 0 180 $X=172820 $Y=454120
X352 982 15 14 983 5 233 984 43 985 SDFFRXL $T=174000 449500 1 0 $X=173400 $Y=443680
X353 986 15 14 987 5 233 988 43 989 SDFFRXL $T=175160 449500 0 0 $X=174560 $Y=449140
X354 990 15 14 991 5 233 992 39 993 SDFFRXL $T=196040 491260 1 180 $X=174560 $Y=490900
X355 994 15 14 995 5 233 996 43 997 SDFFRXL $T=198360 428620 0 0 $X=197760 $Y=428260
X356 998 15 14 999 5 233 1000 43 1001 SDFFRXL $T=198360 439060 0 0 $X=197760 $Y=438700
X357 1002 15 14 1003 5 233 1004 43 1005 SDFFRXL $T=198360 449500 0 0 $X=197760 $Y=449140
X358 1006 15 14 1007 5 233 1008 39 1009 SDFFRXL $T=198360 491260 0 0 $X=197760 $Y=490900
X359 1010 15 14 1011 5 233 1012 39 1013 SDFFRXL $T=198360 501700 1 0 $X=197760 $Y=495880
X360 1014 15 14 1015 5 233 1016 27 1017 SDFFRXL $T=198360 522580 0 0 $X=197760 $Y=522220
X361 1018 15 14 1019 5 233 1020 27 1021 SDFFRXL $T=198360 533020 1 0 $X=197760 $Y=527200
X362 1022 15 14 1023 5 233 1024 43 1025 SDFFRXL $T=223300 439060 0 180 $X=201820 $Y=433240
X363 1026 15 14 1027 5 233 1028 39 1029 SDFFRXL $T=223300 491260 0 180 $X=201820 $Y=485440
X364 1030 15 14 1031 5 233 1032 43 1033 SDFFRXL $T=208800 407740 0 0 $X=208200 $Y=407380
X365 1034 15 14 93 5 97 1035 45 1035 SDFFRXL $T=234900 397300 0 180 $X=213420 $Y=391480
X366 1036 15 14 1037 5 233 1038 27 1039 SDFFRXL $T=215180 522580 1 0 $X=214580 $Y=516760
X367 1040 15 14 84 5 233 1041 45 1042 SDFFRXL $T=217500 428620 1 0 $X=216900 $Y=422800
X368 1043 15 14 1044 5 233 1045 43 1046 SDFFRXL $T=219240 428620 0 0 $X=218640 $Y=428260
X369 1047 15 14 1048 5 233 1049 27 1050 SDFFRXL $T=219240 522580 0 0 $X=218640 $Y=522220
X370 1051 15 14 1052 5 233 1053 39 1054 SDFFRXL $T=220400 491260 0 0 $X=219800 $Y=490900
X371 94 15 14 95 5 97 1055 45 1056 SDFFRXL $T=222140 386860 1 0 $X=221540 $Y=381040
X372 1057 15 14 96 5 97 1058 45 1059 SDFFRXL $T=222140 386860 0 0 $X=221540 $Y=386500
X373 1060 15 14 80 5 233 1061 43 1062 SDFFRXL $T=222720 439060 0 0 $X=222120 $Y=438700
X374 1063 15 14 1064 5 233 1065 43 1066 SDFFRXL $T=223300 439060 1 0 $X=222700 $Y=433240
X375 1067 15 14 1068 5 233 1069 39 1070 SDFFRXL $T=244180 491260 0 180 $X=222700 $Y=485440
X376 1071 15 14 1072 5 233 1073 27 1074 SDFFRXL $T=229680 512140 0 0 $X=229080 $Y=511780
X377 1075 15 14 1076 5 233 1077 39 1078 SDFFRXL $T=232580 480820 0 0 $X=231980 $Y=480460
X378 1079 15 14 1080 5 233 1081 43 1082 SDFFRXL $T=240120 428620 0 0 $X=239520 $Y=428260
X379 1083 15 14 1084 5 233 1085 27 1086 SDFFRXL $T=240120 522580 0 0 $X=239520 $Y=522220
X380 103 15 14 105 5 97 1087 45 1088 SDFFRXL $T=241860 397300 1 0 $X=241260 $Y=391480
X381 1089 15 14 104 5 97 1090 45 1091 SDFFRXL $T=243020 386860 0 0 $X=242420 $Y=386500
X382 98 15 14 106 5 233 1092 45 1093 SDFFRXL $T=243600 386860 1 0 $X=243000 $Y=381040
X383 1094 15 14 1095 5 233 1096 43 1097 SDFFRXL $T=244180 428620 1 0 $X=243580 $Y=422800
X384 1098 15 14 75 5 233 1099 43 1100 SDFFRXL $T=244180 439060 1 0 $X=243580 $Y=433240
X385 1101 15 14 1102 5 233 1103 39 1104 SDFFRXL $T=244180 491260 1 0 $X=243580 $Y=485440
X386 1105 15 14 1106 5 233 1107 39 1108 SDFFRXL $T=251720 491260 0 0 $X=251120 $Y=490900
X387 1109 15 14 1110 5 233 1111 27 1112 SDFFRXL $T=252300 533020 1 0 $X=251700 $Y=527200
X388 1113 15 14 1114 5 233 1115 39 1116 SDFFRXL $T=253460 480820 0 0 $X=252860 $Y=480460
X389 108 15 14 109 5 97 1117 45 1118 SDFFRXL $T=254040 376420 0 0 $X=253440 $Y=376060
X390 1119 15 14 1120 5 233 1121 27 1122 SDFFRXL $T=255780 522580 1 0 $X=255180 $Y=516760
X391 111 15 14 110 5 97 1123 45 1124 SDFFRXL $T=265060 386860 1 0 $X=264460 $Y=381040
X392 1125 15 14 1126 5 233 1127 43 1128 SDFFRXL $T=265060 428620 1 0 $X=264460 $Y=422800
X393 1129 15 14 1130 5 233 1131 43 1132 SDFFRXL $T=265060 428620 0 0 $X=264460 $Y=428260
X394 1133 15 14 1134 5 233 1135 43 1136 SDFFRXL $T=265060 439060 1 0 $X=264460 $Y=433240
X395 1137 15 14 1138 5 233 1139 39 1140 SDFFRXL $T=265060 491260 1 0 $X=264460 $Y=485440
X396 1141 15 14 1142 5 234 306 313 307 SDFFRXL $T=378160 501700 0 0 $X=377560 $Y=501340
X397 1143 15 14 1144 5 234 329 1145 328 SDFFRXL $T=399040 439060 0 0 $X=398440 $Y=438700
X398 1146 15 14 1147 5 234 319 343 318 SDFFRXL $T=399040 501700 0 0 $X=398440 $Y=501340
X399 1148 15 14 1149 5 234 338 337 339 SDFFRXL $T=400200 439060 1 0 $X=399600 $Y=433240
X400 1150 15 14 1151 5 235 350 1152 351 SDFFRXL $T=421660 501700 0 0 $X=421060 $Y=501340
X401 1153 15 14 1154 5 234 384 365 385 SDFFRXL $T=436740 449500 1 0 $X=436140 $Y=443680
X402 1155 15 14 1156 5 235 380 373 381 SDFFRXL $T=437320 512140 1 0 $X=436720 $Y=506320
X403 75 1030 15 14 237 73 XNOR3X1 $T=178640 376420 1 180 $X=160640 $Y=376060
X404 75 1030 15 14 238 76 XNOR3X1 $T=188500 386860 0 180 $X=170500 $Y=381040
X405 1095 75 15 14 1157 88 XNOR3X1 $T=198360 376420 0 0 $X=197760 $Y=376060
X406 1095 1098 15 14 1158 90 XNOR3X1 $T=204740 386860 1 0 $X=204140 $Y=381040
X407 1105 1026 15 14 243 1032 XNOR3X1 $T=207060 449500 1 0 $X=206460 $Y=443680
X408 1106 1026 15 14 241 1033 XNOR3X1 $T=213440 459940 0 0 $X=212840 $Y=459580
X409 614 618 15 14 1159 1085 XNOR3X1 $T=236060 543460 0 0 $X=235460 $Y=543100
X410 1138 1106 15 14 1160 1096 XNOR3X1 $T=244760 439060 0 0 $X=244160 $Y=438700
X411 1138 1105 15 14 1161 1097 XNOR3X1 $T=249980 459940 0 0 $X=249380 $Y=459580
X412 1106 1137 15 14 1162 1099 XNOR3X1 $T=268540 449500 0 180 $X=250540 $Y=443680
X413 1120 1084 15 14 1163 1107 XNOR3X1 $T=251140 512140 1 0 $X=250540 $Y=506320
X414 75 1095 15 14 1164 1093 XNOR3X1 $T=254620 397300 0 0 $X=254020 $Y=396940
X415 618 614 15 14 1165 1122 XNOR3X1 $T=256940 543460 0 0 $X=256340 $Y=543100
X416 75 1094 15 14 1166 1092 XNOR3X1 $T=259840 407740 1 0 $X=259240 $Y=401920
X417 1095 1129 15 14 249 114 XNOR3X1 $T=265640 397300 1 0 $X=265040 $Y=391480
X418 1095 1129 15 14 250 116 XNOR3X1 $T=266800 386860 0 0 $X=266200 $Y=386500
X419 1106 1138 15 14 1167 1100 XNOR3X1 $T=268540 449500 1 0 $X=267940 $Y=443680
X420 1137 1075 15 14 245 1132 XNOR3X1 $T=268540 470380 0 0 $X=267940 $Y=470020
X421 1138 1075 15 14 247 1131 XNOR3X1 $T=268540 480820 1 0 $X=267940 $Y=475000
X422 1084 1120 15 14 1168 1140 XNOR3X1 $T=268540 512140 1 0 $X=267940 $Y=506320
X423 620 714 15 14 1169 440 XNOR3X1 $T=300440 522580 1 0 $X=299840 $Y=516760
X424 623 555 15 14 1170 439 XNOR3X1 $T=318420 533020 0 180 $X=300420 $Y=527200
X425 636 714 15 14 1171 438 XNOR3X1 $T=319000 533020 1 180 $X=301000 $Y=532660
X426 626 723 15 14 1172 624 XNOR3X1 $T=325380 480820 0 180 $X=307380 $Y=475000
X427 629 723 15 14 1173 621 XNOR3X1 $T=327700 480820 1 180 $X=309700 $Y=480460
X428 632 1174 15 14 1175 640 XNOR3X1 $T=317260 397300 0 0 $X=316660 $Y=396940
X429 645 1174 15 14 1176 627 XNOR3X1 $T=334660 418180 1 180 $X=316660 $Y=417820
X430 634 1174 15 14 1177 630 XNOR3X1 $T=317840 428620 1 0 $X=317240 $Y=422800
X431 639 723 15 14 1178 643 XNOR3X1 $T=320160 459940 1 0 $X=319560 $Y=454120
X432 652 555 15 14 1179 442 XNOR3X1 $T=337560 533020 1 180 $X=319560 $Y=532660
X433 642 714 15 14 1180 443 XNOR3X1 $T=320740 512140 1 0 $X=320140 $Y=506320
X434 658 723 15 14 1181 637 XNOR3X1 $T=339300 491260 0 180 $X=321300 $Y=485440
X435 671 555 15 14 1182 441 XNOR3X1 $T=344520 543460 0 180 $X=326520 $Y=537640
X436 655 723 15 14 1183 650 XNOR3X1 $T=336980 459940 0 0 $X=336380 $Y=459580
X437 649 555 15 14 1184 444 XNOR3X1 $T=338720 512140 1 0 $X=338120 $Y=506320
X438 676 1174 15 14 1185 659 XNOR3X1 $T=339300 418180 0 0 $X=338700 $Y=417820
X439 661 723 15 14 1186 653 XNOR3X1 $T=339880 501700 1 0 $X=339280 $Y=495880
X440 667 555 15 14 1187 445 XNOR3X1 $T=339880 543460 0 0 $X=339280 $Y=543100
X441 647 1174 15 14 1188 656 XNOR3X1 $T=341040 407740 1 0 $X=340440 $Y=401920
X442 678 1174 15 14 1189 662 XNOR3X1 $T=351480 428620 0 0 $X=350880 $Y=428260
X443 664 723 15 14 1190 668 XNOR3X1 $T=354380 459940 0 0 $X=353780 $Y=459580
X444 701 723 15 14 1191 672 XNOR3X1 $T=354960 491260 0 0 $X=354360 $Y=490900
X445 674 716 15 14 1192 665 XNOR3X1 $T=358440 397300 1 0 $X=357840 $Y=391480
X446 686 723 15 14 1193 681 XNOR3X1 $T=375840 501700 0 180 $X=357840 $Y=495880
X447 699 1174 15 14 1194 687 XNOR3X1 $T=378160 428620 0 0 $X=377560 $Y=428260
X448 703 723 15 14 1195 690 XNOR3X1 $T=378160 491260 0 0 $X=377560 $Y=490900
X449 1142 714 15 14 1196 447 XNOR3X1 $T=378160 543460 1 0 $X=377560 $Y=537640
X450 694 1174 15 14 1197 702 XNOR3X1 $T=378740 439060 1 0 $X=378140 $Y=433240
X451 696 714 15 14 1198 446 XNOR3X1 $T=379900 533020 0 0 $X=379300 $Y=532660
X452 709 1174 15 14 1199 705 XNOR3X1 $T=395560 428620 0 0 $X=394960 $Y=428260
X453 712 555 15 14 1200 448 XNOR3X1 $T=413540 543460 0 180 $X=395540 $Y=537640
X454 1147 714 15 14 1201 449 XNOR3X1 $T=401940 522580 1 0 $X=401340 $Y=516760
X455 744 723 15 14 1202 713 XNOR3X1 $T=424560 501700 0 180 $X=406560 $Y=495880
X456 726 564 15 14 1203 450 XNOR3X1 $T=419920 543460 1 0 $X=419320 $Y=537640
X457 734 731 15 14 1204 727 XNOR3X1 $T=421660 491260 0 0 $X=421060 $Y=490900
X458 717 158 15 14 1205 735 XNOR3X1 $T=424560 439060 1 0 $X=423960 $Y=433240
X459 162 1174 15 14 1206 745 XNOR3X1 $T=436160 407740 1 0 $X=435560 $Y=401920
X460 1156 728 15 14 1207 452 XNOR3X1 $T=437320 543460 1 0 $X=436720 $Y=537640
X461 461 728 15 14 1208 454 XNOR3X1 $T=465740 533020 1 180 $X=447740 $Y=532660
X462 759 158 15 14 1209 763 XNOR3X1 $T=468060 428620 0 0 $X=467460 $Y=428260
X463 458 730 15 14 1210 456 XNOR3X1 $T=468060 459940 0 0 $X=467460 $Y=459580
X464 762 730 15 14 1211 766 XNOR3X1 $T=468060 491260 0 0 $X=467460 $Y=490900
X465 175 160 15 14 1212 459 XNOR3X1 $T=470380 397300 1 0 $X=469780 $Y=391480
X466 765 728 15 14 1213 457 XNOR3X1 $T=470380 533020 0 0 $X=469780 $Y=532660
X467 779 731 15 14 1214 769 XNOR3X1 $T=473860 501700 1 0 $X=473260 $Y=495880
X468 183 158 15 14 179 775 XNOR3X1 $T=499380 386860 0 180 $X=481380 $Y=381040
X469 777 158 15 14 1215 780 XNOR3X1 $T=485460 428620 0 0 $X=484860 $Y=428260
X470 782 1216 15 14 1217 772 XNOR3X1 $T=487200 428620 1 0 $X=486600 $Y=422800
X471 784 564 15 14 1218 463 XNOR3X1 $T=487780 533020 0 0 $X=487180 $Y=532660
X472 787 728 15 14 1219 464 XNOR3X1 $T=489520 543460 0 0 $X=488920 $Y=543100
X473 771 730 15 14 1220 785 XNOR3X1 $T=490100 491260 0 0 $X=489500 $Y=490900
X474 792 731 15 14 1221 788 XNOR3X1 $T=494160 501700 1 0 $X=493560 $Y=495880
X475 774 731 15 14 1222 462 XNOR3X1 $T=514460 449500 1 180 $X=496460 $Y=449140
X476 806 728 15 14 421 465 XNOR3X1 $T=502280 543460 1 0 $X=501680 $Y=537640
X477 790 158 15 14 1223 793 XNOR3X1 $T=502860 428620 0 0 $X=502260 $Y=428260
X478 795 728 15 14 1224 466 XNOR3X1 $T=505180 533020 0 0 $X=504580 $Y=532660
X479 799 731 15 14 1225 796 XNOR3X1 $T=507500 491260 0 0 $X=506900 $Y=490900
X480 191 158 15 14 1226 801 XNOR3X1 $T=509240 428620 1 0 $X=508640 $Y=422800
X481 818 731 15 14 1227 810 XNOR3X1 $T=522000 501700 1 0 $X=521400 $Y=495880
X482 202 158 15 14 1228 816 XNOR3X1 $T=522580 418180 1 0 $X=521980 $Y=412360
X483 803 731 15 14 1229 813 XNOR3X1 $T=522580 449500 1 0 $X=521980 $Y=443680
X484 809 564 15 14 1230 468 XNOR3X1 $T=522580 543460 1 0 $X=521980 $Y=537640
X485 198 158 15 14 1231 804 XNOR3X1 $T=523160 386860 1 0 $X=522560 $Y=381040
X486 812 564 15 14 1232 467 XNOR3X1 $T=523160 533020 0 0 $X=522560 $Y=532660
X487 815 731 15 14 1233 807 XNOR3X1 $T=524900 491260 0 0 $X=524300 $Y=490900
X488 199 158 15 14 1234 819 XNOR3X1 $T=528380 407740 0 0 $X=527780 $Y=407380
X489 652 15 14 1235 1236 1182 651 555 OAI221XL $T=338140 533020 0 180 $X=331740 $Y=527200
X490 631 15 14 1237 272 1238 1239 269 OAI221XL $T=335820 397300 0 0 $X=335220 $Y=396940
X491 667 15 14 266 265 1184 666 555 OAI221XL $T=346260 522580 1 0 $X=345660 $Y=516760
X492 660 15 14 722 1240 1241 1242 1243 OAI221XL $T=355540 480820 1 0 $X=354940 $Y=475000
X493 677 15 14 1237 1244 1245 1246 1247 OAI221XL $T=366560 407740 0 0 $X=365960 $Y=407380
X494 712 15 14 327 320 558 711 555 OAI221XL $T=408320 533020 1 0 $X=407720 $Y=527200
X495 797 15 14 357 1248 1249 725 1250 OAI221XL $T=435580 522580 1 180 $X=429180 $Y=522220
X496 739 15 14 1251 1248 1207 738 1252 OAI221XL $T=442540 533020 0 0 $X=441940 $Y=532660
X497 768 15 14 1251 1248 1213 767 1253 OAI221XL $T=486620 533020 0 180 $X=480220 $Y=527200
X498 1254 15 14 1255 1216 1256 789 1257 OAI221XL $T=501120 407740 1 0 $X=500520 $Y=401920
X499 806 15 14 1251 1248 1224 805 422 OAI221XL $T=502860 533020 1 0 $X=502260 $Y=527200
X500 1258 15 14 413 1216 1259 194 418 OAI221XL $T=512720 386860 1 0 $X=512120 $Y=381040
X501 1260 15 14 423 730 1261 802 428 OAI221XL $T=516200 449500 0 0 $X=515600 $Y=449140
X502 811 15 14 1262 1263 1230 812 564 OAI221XL $T=533020 522580 1 180 $X=526620 $Y=522220
X503 264 267 15 14 714 1187 OR3X1 $T=346260 522580 0 0 $X=345660 $Y=522220
X504 1264 278 15 14 1265 1266 OR3X1 $T=371200 533020 1 0 $X=370600 $Y=527200
X505 310 797 15 14 1146 320 OR3X1 $T=399620 533020 1 0 $X=399020 $Y=527200
X506 321 326 15 14 714 1200 OR3X1 $T=406000 533020 1 180 $X=400760 $Y=532660
X507 1267 314 15 14 1268 1269 OR3X1 $T=413540 459940 0 0 $X=412940 $Y=459580
X508 1270 1271 15 14 1272 1273 OR3X1 $T=426880 407740 1 0 $X=426280 $Y=401920
X509 1274 1275 15 14 1276 1277 OR3X1 $T=433840 480820 0 180 $X=428600 $Y=475000
X510 1278 1279 15 14 1280 1281 OR3X1 $T=439640 418180 1 180 $X=434400 $Y=417820
X511 1282 420 15 14 408 1283 OR3X1 $T=505760 480820 0 180 $X=500520 $Y=475000
X512 1284 436 15 14 433 1285 OR3X1 $T=522580 418180 0 180 $X=517340 $Y=412360
X513 703 15 14 1286 722 301 1287 OAI211XL $T=386280 480820 0 0 $X=385680 $Y=480460
X514 709 15 14 1288 1237 309 1289 OAI211XL $T=392660 418180 0 0 $X=392060 $Y=417820
X515 723 15 14 1290 1143 315 1291 OAI211XL $T=401940 459940 0 0 $X=401340 $Y=459580
X516 361 15 14 559 1248 1292 1293 OAI211XL $T=444860 533020 0 180 $X=440200 $Y=527200
X517 759 15 14 1294 1216 1295 1296 OAI211XL $T=468060 418180 0 0 $X=467460 $Y=417820
X518 761 15 14 1297 730 1298 1299 OAI211XL $T=468060 480820 0 0 $X=467460 $Y=480460
X519 679 15 14 798 714 1300 279 797 OAI32XL $T=360760 533020 1 0 $X=360160 $Y=527200
X520 1301 15 14 333 335 338 1302 135 OAI32XL $T=412960 418180 0 0 $X=412360 $Y=417820
X521 798 15 14 1303 1304 1203 356 797 OAI32XL $T=428040 533020 1 0 $X=427440 $Y=527200
X522 1305 15 14 371 367 1152 1306 125 OAI32XL $T=441380 491260 1 0 $X=440780 $Y=485440
X523 1307 15 14 383 379 376 1308 126 OAI32XL $T=455300 428620 0 180 $X=449480 $Y=422800
X524 1309 15 14 1310 1311 OR2X1 $T=175160 386860 0 0 $X=174560 $Y=386500
X525 1312 15 14 1313 79 OR2X1 $T=192560 386860 0 180 $X=188480 $Y=381040
X526 1098 15 14 1030 1314 OR2X1 $T=201840 397300 0 180 $X=197760 $Y=391480
X527 75 15 14 80 1315 OR2X1 $T=201260 386860 0 0 $X=200660 $Y=386500
X528 1105 15 14 1026 1316 OR2X1 $T=213440 459940 1 0 $X=212840 $Y=454120
X529 1040 15 14 93 1317 OR2X1 $T=218080 386860 0 0 $X=217480 $Y=386500
X530 1318 15 14 1319 1320 OR2X1 $T=220400 470380 0 0 $X=219800 $Y=470020
X531 1321 15 14 1322 1323 OR2X1 $T=243600 449500 1 180 $X=239520 $Y=449140
X532 1106 15 14 1068 1324 OR2X1 $T=254620 459940 0 180 $X=250540 $Y=454120
X533 1325 15 14 1326 1327 OR2X1 $T=263320 470380 1 0 $X=262720 $Y=464560
X534 1138 15 14 1114 1328 OR2X1 $T=276660 459940 1 0 $X=276060 $Y=454120
X535 1329 15 14 1330 1331 OR2X1 $T=284780 459940 0 180 $X=280700 $Y=454120
X536 1332 15 14 1333 1334 OR2X1 $T=291740 418180 0 180 $X=287660 $Y=412360
X537 1137 15 14 1075 1335 OR2X1 $T=289420 470380 0 0 $X=288820 $Y=470020
X538 1094 15 14 1129 1336 OR2X1 $T=291160 407740 1 0 $X=290560 $Y=401920
X539 1337 15 14 1338 1339 OR2X1 $T=305080 386860 1 180 $X=301000 $Y=386500
X540 1095 15 14 1126 1340 OR2X1 $T=305660 397300 0 180 $X=301580 $Y=391480
X541 1341 15 14 1342 1170 OR2X1 $T=310300 522580 1 180 $X=306220 $Y=522220
X542 628 15 14 625 1343 OR2X1 $T=316680 459940 1 0 $X=316080 $Y=454120
X543 723 15 14 629 1344 OR2X1 $T=317840 470380 1 0 $X=317240 $Y=464560
X544 1174 15 14 634 1345 OR2X1 $T=322480 418180 1 0 $X=321880 $Y=412360
X545 255 15 14 1346 1347 OR2X1 $T=326540 522580 0 180 $X=322460 $Y=516760
X546 629 15 14 626 1348 OR2X1 $T=325380 480820 1 0 $X=324780 $Y=475000
X547 633 15 14 644 1349 OR2X1 $T=327120 397300 1 0 $X=326520 $Y=391480
X548 1347 15 14 1350 1351 OR2X1 $T=327120 522580 1 0 $X=326520 $Y=516760
X549 723 15 14 639 1352 OR2X1 $T=327700 449500 0 0 $X=327100 $Y=449140
X550 1353 15 14 798 1235 OR2X1 $T=327700 522580 0 0 $X=327100 $Y=522220
X551 634 15 14 645 1354 OR2X1 $T=331180 407740 0 0 $X=330580 $Y=407380
X552 1351 15 14 797 1236 OR2X1 $T=331760 522580 0 0 $X=331160 $Y=522220
X553 1353 15 14 1355 1356 OR2X1 $T=335820 522580 0 0 $X=335220 $Y=522220
X554 723 15 14 654 1357 OR2X1 $T=341620 449500 0 180 $X=337540 $Y=443680
X555 646 15 14 1174 1358 OR2X1 $T=343360 397300 0 180 $X=339280 $Y=391480
X556 1359 15 14 1360 1186 OR2X1 $T=343360 480820 0 0 $X=342760 $Y=480460
X557 722 15 14 657 1243 OR2X1 $T=353800 480820 0 180 $X=349720 $Y=475000
X558 723 15 14 657 1361 OR2X1 $T=357280 491260 0 180 $X=353200 $Y=485440
X559 798 15 14 553 266 OR2X1 $T=357860 522580 1 180 $X=353780 $Y=522220
X560 1237 15 14 675 1247 OR2X1 $T=357860 407740 0 0 $X=357260 $Y=407380
X561 1351 15 14 1362 1264 OR2X1 $T=357860 522580 0 0 $X=357260 $Y=522220
X562 1174 15 14 675 1363 OR2X1 $T=359600 418180 1 0 $X=359000 $Y=412360
X563 556 15 14 1300 557 OR2X1 $T=363660 543460 1 0 $X=363060 $Y=537640
X564 1364 15 14 1365 1189 OR2X1 $T=367720 418180 0 180 $X=363640 $Y=412360
X565 700 15 14 685 1366 OR2X1 $T=375840 470380 1 180 $X=371760 $Y=470020
X566 723 15 14 701 1367 OR2X1 $T=382220 491260 0 180 $X=378140 $Y=485440
X567 701 15 14 686 1368 OR2X1 $T=379320 470380 1 0 $X=378720 $Y=464560
X568 1174 15 14 694 1369 OR2X1 $T=379900 428620 1 0 $X=379300 $Y=422800
X569 1356 15 14 1370 1371 OR2X1 $T=379900 522580 0 0 $X=379300 $Y=522220
X570 736 15 14 692 1372 OR2X1 $T=383960 386860 1 180 $X=379880 $Y=386500
X571 693 15 14 698 296 OR2X1 $T=385120 407740 0 180 $X=381040 $Y=401920
X572 736 15 14 691 1373 OR2X1 $T=387440 386860 0 180 $X=383360 $Y=381040
X573 694 15 14 699 1374 OR2X1 $T=387440 407740 1 0 $X=386840 $Y=401920
X574 1266 15 14 1375 310 OR2X1 $T=392660 533020 1 0 $X=392060 $Y=527200
X575 1376 15 14 1377 306 OR2X1 $T=400780 480820 0 180 $X=396700 $Y=475000
X576 707 15 14 704 1378 OR2X1 $T=401940 459940 0 180 $X=397860 $Y=454120
X577 706 15 14 1143 1379 OR2X1 $T=400200 470380 0 0 $X=399600 $Y=470020
X578 1144 15 14 1149 1380 OR2X1 $T=404260 459940 1 0 $X=403660 $Y=454120
X579 710 15 14 719 1381 OR2X1 $T=406000 397300 1 0 $X=405400 $Y=391480
X580 1382 15 14 1383 1145 OR2X1 $T=408320 418180 1 0 $X=407720 $Y=412360
X581 755 15 14 721 1384 OR2X1 $T=424560 397300 0 180 $X=420480 $Y=391480
X582 723 15 14 744 1385 OR2X1 $T=421080 470380 0 0 $X=420480 $Y=470020
X583 158 15 14 717 1386 OR2X1 $T=425140 428620 1 0 $X=424540 $Y=422800
X584 731 15 14 734 1387 OR2X1 $T=429200 491260 1 0 $X=428600 $Y=485440
X585 739 15 14 1156 360 OR2X1 $T=440800 522580 1 180 $X=436720 $Y=522220
X586 560 15 14 1154 1388 OR2X1 $T=442540 480820 0 180 $X=438460 $Y=475000
X587 1174 15 14 162 1389 OR2X1 $T=443120 407740 1 180 $X=439040 $Y=407380
X588 737 15 14 742 1390 OR2X1 $T=446020 407740 0 0 $X=445420 $Y=407380
X589 1391 15 14 797 1292 OR2X1 $T=452980 522580 1 180 $X=448900 $Y=522220
X590 749 15 14 1153 1392 OR2X1 $T=455300 470380 1 180 $X=451220 $Y=470020
X591 1393 15 14 1394 380 OR2X1 $T=458200 491260 1 180 $X=454120 $Y=490900
X592 741 15 14 756 1395 OR2X1 $T=455880 407740 1 0 $X=455280 $Y=401920
X593 1396 15 14 1397 384 OR2X1 $T=461100 428620 1 180 $X=457020 $Y=428260
X594 743 15 14 747 1398 OR2X1 $T=457620 459940 1 0 $X=457020 $Y=454120
X595 762 15 14 750 1399 OR2X1 $T=460520 470380 0 0 $X=459920 $Y=470020
X596 743 15 14 746 396 OR2X1 $T=461680 459940 1 0 $X=461080 $Y=454120
X597 760 15 14 757 1400 OR2X1 $T=471540 418180 0 180 $X=467460 $Y=412360
X598 728 15 14 798 1251 OR2X1 $T=468060 533020 1 0 $X=467460 $Y=527200
X599 754 15 14 753 176 OR2X1 $T=470380 386860 0 0 $X=469780 $Y=386500
X600 392 15 14 1401 1402 OR2X1 $T=475020 522580 0 0 $X=474420 $Y=522220
X601 770 15 14 778 402 OR2X1 $T=483720 480820 1 0 $X=483120 $Y=475000
X602 782 15 14 777 1403 OR2X1 $T=485460 418180 0 0 $X=484860 $Y=417820
X603 771 15 14 779 1404 OR2X1 $T=488940 491260 1 180 $X=484860 $Y=490900
X604 781 15 14 776 404 OR2X1 $T=488360 397300 1 0 $X=487760 $Y=391480
X605 410 15 14 1405 1406 OR2X1 $T=493580 522580 1 180 $X=489500 $Y=522220
X606 728 15 14 797 1248 OR2X1 $T=490100 533020 1 0 $X=489500 $Y=527200
X607 1407 15 14 728 1218 OR2X1 $T=496480 533020 1 0 $X=495880 $Y=527200
X608 412 15 14 1408 1409 OR2X1 $T=502280 522580 0 180 $X=498200 $Y=516760
X609 731 15 14 799 407 OR2X1 $T=504020 480820 0 0 $X=503420 $Y=480460
X610 1216 15 14 189 1257 OR2X1 $T=505180 397300 0 0 $X=504580 $Y=396940
X611 1410 15 14 1411 1221 OR2X1 $T=505180 491260 1 0 $X=504580 $Y=485440
X612 1412 15 14 1413 1223 OR2X1 $T=506920 407740 1 0 $X=506320 $Y=401920
X613 773 15 14 731 1414 OR2X1 $T=506920 439060 0 0 $X=506320 $Y=438700
X614 1415 15 14 731 419 OR2X1 $T=516780 480820 0 180 $X=512700 $Y=475000
X615 1416 15 14 1417 1418 OR2X1 $T=517360 522580 0 180 $X=513280 $Y=516760
X616 1402 15 14 797 1263 OR2X1 $T=516200 522580 0 0 $X=515600 $Y=522220
X617 1402 15 14 1419 1420 OR2X1 $T=518520 533020 1 0 $X=517920 $Y=527200
X618 1415 15 14 730 1421 OR2X1 $T=522580 470380 1 180 $X=518500 $Y=470020
X619 1416 15 14 798 1262 OR2X1 $T=520840 522580 0 0 $X=520240 $Y=522220
X620 158 15 14 199 1422 OR2X1 $T=522000 397300 0 0 $X=521400 $Y=396940
X621 199 15 14 202 1423 OR2X1 $T=526060 407740 0 180 $X=521980 $Y=401920
X622 817 15 14 814 1424 OR2X1 $T=528960 459940 1 180 $X=524880 $Y=459580
X623 731 15 14 818 1425 OR2X1 $T=527220 491260 1 0 $X=526620 $Y=485440
X624 1426 1427 15 14 1309 NOR2BXL $T=171680 386860 0 0 $X=171080 $Y=386500
X625 1427 75 15 14 1031 NOR2BXL $T=175740 397300 1 0 $X=175140 $Y=391480
X626 1428 1031 15 14 1098 NOR2BXL $T=191980 397300 1 0 $X=191380 $Y=391480
X627 1429 1098 15 14 80 NOR2BXL $T=196040 386860 0 180 $X=191960 $Y=381040
X628 1430 1431 15 14 1311 NOR2BXL $T=192560 386860 0 0 $X=191960 $Y=386500
X629 1312 239 15 14 1432 NOR2BXL $T=201840 397300 1 0 $X=201240 $Y=391480
X630 1433 75 15 14 80 NOR2BXL $T=208800 397300 0 0 $X=208200 $Y=396940
X631 1434 1435 15 14 1318 NOR2BXL $T=219820 480820 0 180 $X=215740 $Y=475000
X632 1436 1027 15 14 1105 NOR2BXL $T=222720 459940 0 180 $X=218640 $Y=454120
X633 1435 1106 15 14 1027 NOR2BXL $T=220400 480820 1 0 $X=219800 $Y=475000
X634 1321 243 15 14 1437 NOR2BXL $T=237220 449500 1 180 $X=233140 $Y=449140
X635 1438 1439 15 14 1320 NOR2BXL $T=239540 459940 1 180 $X=235460 $Y=459580
X636 1440 1106 15 14 1068 NOR2BXL $T=249400 470380 0 180 $X=245320 $Y=464560
X637 1441 1105 15 14 1068 NOR2BXL $T=250560 449500 0 0 $X=249960 $Y=449140
X638 1442 1138 15 14 1076 NOR2BXL $T=262160 470380 1 180 $X=258080 $Y=470020
X639 1443 1442 15 14 1325 NOR2BXL $T=266800 470380 1 180 $X=262720 $Y=470020
X640 1444 1138 15 14 1114 NOR2BXL $T=268540 449500 1 180 $X=264460 $Y=449140
X641 1445 1446 15 14 1327 NOR2BXL $T=275500 459940 0 180 $X=271420 $Y=454120
X642 1447 1095 15 14 1126 NOR2BXL $T=273760 418180 1 0 $X=273160 $Y=412360
X643 1448 1137 15 14 1114 NOR2BXL $T=278400 459940 1 180 $X=274320 $Y=459580
X644 1329 245 15 14 1449 NOR2BXL $T=285360 470380 0 180 $X=281280 $Y=464560
X645 1450 1451 15 14 1334 NOR2BXL $T=291740 407740 1 180 $X=287660 $Y=407380
X646 1452 1076 15 14 1137 NOR2BXL $T=292320 470380 0 180 $X=288240 $Y=464560
X647 1337 251 15 14 1453 NOR2BXL $T=299860 397300 1 180 $X=295780 $Y=396940
X648 1454 1130 15 14 1094 NOR2BXL $T=296960 418180 1 0 $X=296360 $Y=412360
X649 1455 1094 15 14 1126 NOR2BXL $T=303920 407740 0 180 $X=299840 $Y=401920
X650 1456 1457 15 14 1332 NOR2BXL $T=304500 418180 0 180 $X=300420 $Y=412360
X651 1457 1095 15 14 1130 NOR2BXL $T=302180 407740 0 0 $X=301580 $Y=407380
X652 1169 1458 15 14 555 NOR2BXL $T=314940 512140 0 0 $X=314340 $Y=511780
X653 1341 1347 15 14 798 NOR2BXL $T=318420 522580 1 0 $X=317820 $Y=516760
X654 1342 798 15 14 1459 NOR2BXL $T=319000 522580 0 0 $X=318400 $Y=522220
X655 1459 256 15 14 1460 NOR2BXL $T=323060 512140 1 180 $X=318980 $Y=511780
X656 260 722 15 14 1348 NOR2BXL $T=333500 480820 0 180 $X=329420 $Y=475000
X657 1461 1462 15 14 1357 NOR2BXL $T=335240 449500 0 180 $X=331160 $Y=443680
X658 1239 1174 15 14 631 NOR2BXL $T=335820 397300 0 180 $X=331740 $Y=391480
X659 1463 1464 15 14 1358 NOR2BXL $T=336400 397300 1 0 $X=335800 $Y=391480
X660 270 1237 15 14 1354 NOR2BXL $T=344520 407740 1 180 $X=340440 $Y=407380
X661 268 1237 15 14 647 NOR2BXL $T=345100 397300 1 180 $X=341020 $Y=396940
X662 1465 722 15 14 655 NOR2BXL $T=343940 459940 1 0 $X=343340 $Y=454120
X663 264 797 15 14 553 NOR2BXL $T=350900 522580 0 0 $X=350300 $Y=522220
X664 1242 723 15 14 660 NOR2BXL $T=361340 470380 0 0 $X=360740 $Y=470020
X665 282 1241 15 14 261 NOR2BXL $T=367140 480820 0 180 $X=363060 $Y=475000
X666 288 1245 15 14 271 NOR2BXL $T=371200 418180 0 180 $X=367120 $Y=412360
X667 278 714 15 14 679 NOR2BXL $T=367720 533020 1 0 $X=367120 $Y=527200
X668 280 683 15 14 734 NOR2BXL $T=369460 459940 1 0 $X=368860 $Y=454120
X669 1246 1174 15 14 677 NOR2BXL $T=372360 407740 0 0 $X=371760 $Y=407380
X670 290 733 15 14 683 NOR2BXL $T=378160 459940 1 0 $X=377560 $Y=454120
X671 1466 723 15 14 1368 NOR2BXL $T=386280 470380 0 180 $X=382200 $Y=464560
X672 1196 1467 15 14 555 NOR2BXL $T=387440 533020 1 0 $X=386840 $Y=527200
X673 1468 1371 15 14 1469 NOR2BXL $T=393820 522580 1 180 $X=389740 $Y=522220
X674 300 722 15 14 1368 NOR2BXL $T=394980 470380 1 180 $X=390900 $Y=470020
X675 308 1237 15 14 1374 NOR2BXL $T=396140 407740 0 180 $X=392060 $Y=401920
X676 1470 1174 15 14 1374 NOR2BXL $T=404260 407740 0 180 $X=400180 $Y=401920
X677 1471 722 15 14 1380 NOR2BXL $T=411220 470380 0 180 $X=407140 $Y=464560
X678 344 720 15 14 719 NOR2BXL $T=414120 397300 0 180 $X=410040 $Y=391480
X679 1268 723 15 14 1380 NOR2BXL $T=421660 459940 1 180 $X=417580 $Y=459580
X680 1472 1237 15 14 1384 NOR2BXL $T=419920 407740 1 0 $X=419320 $Y=401920
X681 1272 1174 15 14 1384 NOR2BXL $T=426880 407740 0 180 $X=422800 $Y=401920
X682 1276 731 15 14 1388 NOR2BXL $T=431520 480820 0 0 $X=430920 $Y=480460
X683 1473 730 15 14 1388 NOR2BXL $T=439060 480820 0 0 $X=438460 $Y=480460
X684 1474 1216 15 14 1390 NOR2BXL $T=444860 418180 0 0 $X=444260 $Y=417820
X685 1280 158 15 14 1390 NOR2BXL $T=445440 418180 1 0 $X=444840 $Y=412360
X686 370 1475 15 14 125 NOR2BXL $T=456460 491260 1 0 $X=455860 $Y=485440
X687 382 1476 15 14 126 NOR2BXL $T=462260 428620 1 0 $X=461660 $Y=422800
X688 398 754 15 14 753 NOR2BXL $T=474440 386860 0 180 $X=470360 $Y=381040
X689 1477 731 15 14 1404 NOR2BXL $T=470960 491260 1 0 $X=470360 $Y=485440
X690 392 728 15 14 455 NOR2BXL $T=471540 522580 0 0 $X=470940 $Y=522220
X691 1478 1409 15 14 1479 NOR2BXL $T=478500 522580 0 0 $X=477900 $Y=522220
X692 1391 1406 15 14 1480 NOR2BXL $T=481980 522580 0 0 $X=481380 $Y=522220
X693 1481 158 15 14 1403 NOR2BXL $T=488940 418180 0 0 $X=488340 $Y=417820
X694 417 1216 15 14 183 NOR2BXL $T=504020 386860 0 180 $X=499940 $Y=381040
X695 1254 158 15 14 789 NOR2BXL $T=501700 397300 0 0 $X=501100 $Y=396940
X696 1482 1256 15 14 426 NOR2BXL $T=502860 407740 0 0 $X=502260 $Y=407380
X697 427 730 15 14 774 NOR2BXL $T=510400 449500 0 180 $X=506320 $Y=443680
X698 411 1418 15 14 1483 NOR2BXL $T=508660 522580 0 0 $X=508060 $Y=522220
X699 415 730 15 14 800 NOR2BXL $T=509240 470380 1 0 $X=508640 $Y=464560
X700 409 1420 15 14 1484 NOR2BXL $T=512720 522580 0 0 $X=512120 $Y=522220
X701 433 158 15 14 191 NOR2BXL $T=517940 418180 0 180 $X=513860 $Y=412360
X702 1260 731 15 14 802 NOR2BXL $T=516780 449500 1 0 $X=516180 $Y=443680
X703 1485 1486 15 14 1414 NOR2BXL $T=521420 439060 1 180 $X=517340 $Y=438700
X704 1258 158 15 14 194 NOR2BXL $T=519680 386860 1 0 $X=519080 $Y=381040
X705 425 1216 15 14 1423 NOR2BXL $T=521420 407740 0 0 $X=520820 $Y=407380
X706 1415 815 15 14 817 NOR2BXL $T=524900 470380 0 0 $X=524300 $Y=470020
X707 1428 239 15 14 1314 1487 OA21X1 $T=192560 386860 1 180 $X=186740 $Y=386500
X708 1044 1031 15 14 1098 1431 OA21X1 $T=207640 397300 1 0 $X=207040 $Y=391480
X709 1436 243 15 14 1316 1488 OA21X1 $T=222720 459940 1 0 $X=222120 $Y=454120
X710 1052 1027 15 14 1105 1439 OA21X1 $T=230840 459940 0 0 $X=230240 $Y=459580
X711 1102 1076 15 14 1137 1446 OA21X1 $T=268540 459940 0 0 $X=267940 $Y=459580
X712 1134 1130 15 14 1094 1451 OA21X1 $T=275500 407740 0 0 $X=274900 $Y=407380
X713 1454 251 15 14 1336 1489 OA21X1 $T=288840 397300 0 0 $X=288240 $Y=396940
X714 1452 245 15 14 1335 1490 OA21X1 $T=291740 459940 0 0 $X=291140 $Y=459580
X715 619 641 15 14 555 1346 OA21X1 $T=307980 512140 1 0 $X=307380 $Y=506320
X716 635 622 15 14 555 1350 OA21X1 $T=314940 512140 1 0 $X=314340 $Y=506320
X717 636 623 15 14 555 1491 OA21X1 $T=320740 533020 1 0 $X=320140 $Y=527200
X718 671 652 15 14 555 1355 OA21X1 $T=344520 522580 1 180 $X=338700 $Y=522220
X719 655 723 15 14 1492 1493 OA21X1 $T=353220 459940 0 180 $X=347400 $Y=454120
X720 651 670 15 14 555 1362 OA21X1 $T=353800 522580 1 0 $X=353200 $Y=516760
X721 680 689 15 14 555 1370 OA21X1 $T=379900 522580 1 0 $X=379300 $Y=516760
X722 1237 297 15 14 295 1494 OA21X1 $T=385120 407740 0 0 $X=384520 $Y=407380
X723 707 722 15 14 299 1495 OA21X1 $T=392080 470380 1 0 $X=391480 $Y=464560
X724 1496 1287 15 14 322 1377 OA21X1 $T=392080 480820 1 0 $X=391480 $Y=475000
X725 695 1141 15 14 555 1375 OA21X1 $T=392080 522580 1 0 $X=391480 $Y=516760
X726 314 1495 15 14 125 1376 OA21X1 $T=397300 470380 1 0 $X=396700 $Y=464560
X727 710 1237 15 14 1494 1497 OA21X1 $T=399040 397300 1 0 $X=398440 $Y=391480
X728 1498 1289 15 14 332 1383 OA21X1 $T=405420 407740 0 0 $X=404820 $Y=407380
X729 719 1237 15 14 1497 1499 OA21X1 $T=409480 397300 0 0 $X=408880 $Y=396940
X730 1271 1499 15 14 126 1382 OA21X1 $T=414700 407740 0 180 $X=408880 $Y=401920
X731 743 722 15 14 1500 1501 OA21X1 $T=419920 470380 1 180 $X=414100 $Y=470020
X732 1237 344 15 14 1497 1502 OA21X1 $T=415280 397300 1 0 $X=414680 $Y=391480
X733 716 1216 15 14 1503 1504 OA21X1 $T=419920 428620 1 0 $X=419320 $Y=422800
X734 160 1237 15 14 1505 1506 OA21X1 $T=429200 407740 1 180 $X=423380 $Y=407380
X735 755 1237 15 14 1502 352 OA21X1 $T=425720 397300 1 0 $X=425120 $Y=391480
X736 733 730 15 14 1507 1508 OA21X1 $T=431520 480820 1 180 $X=425700 $Y=480460
X737 1151 360 15 14 564 1509 OA21X1 $T=436160 522580 1 0 $X=435560 $Y=516760
X738 1155 738 15 14 564 1510 OA21X1 $T=441380 522580 1 0 $X=440780 $Y=516760
X739 798 1478 15 14 1292 1252 OA21X1 $T=445440 533020 1 0 $X=444840 $Y=527200
X740 1511 1299 15 14 370 1394 OA21X1 $T=451240 491260 1 0 $X=450640 $Y=485440
X741 1275 1512 15 14 129 1393 OA21X1 $T=453560 480820 1 0 $X=452960 $Y=475000
X742 1513 1296 15 14 382 1397 OA21X1 $T=457040 428620 1 0 $X=456440 $Y=422800
X743 750 730 15 14 391 1512 OA21X1 $T=464000 480820 0 180 $X=458180 $Y=475000
X744 757 1216 15 14 1514 1515 OA21X1 $T=459360 418180 1 0 $X=458760 $Y=412360
X745 1279 1515 15 14 135 1396 OA21X1 $T=465740 418180 1 180 $X=459920 $Y=417820
X746 461 562 15 14 564 1401 OA21X1 $T=472700 533020 1 0 $X=472100 $Y=527200
X747 760 1216 15 14 1516 1514 OA21X1 $T=480820 418180 0 180 $X=475000 $Y=412360
X748 784 787 15 14 564 1405 OA21X1 $T=487780 522580 1 0 $X=487180 $Y=516760
X749 1216 405 15 14 1285 1516 OA21X1 $T=493580 407740 1 180 $X=487760 $Y=407380
X750 730 403 15 14 1283 1517 OA21X1 $T=491260 480820 0 0 $X=490660 $Y=480460
X751 783 786 15 14 564 1408 OA21X1 $T=493000 522580 1 0 $X=492400 $Y=516760
X752 808 811 15 14 564 1417 OA21X1 $T=523160 522580 0 180 $X=517340 $Y=516760
X753 809 812 15 14 564 1419 OA21X1 $T=528960 533020 0 180 $X=523140 $Y=527200
X754 798 642 15 14 256 255 1458 797 641 OAI33XL $T=325960 512140 0 0 $X=325360 $Y=511780
X755 798 696 15 14 1371 1266 1467 797 695 OAI33XL $T=383960 522580 0 0 $X=383360 $Y=522220
X756 786 798 15 14 412 410 1407 797 787 OAI33XL $T=494160 522580 0 0 $X=493560 $Y=522220
X757 253 1173 15 14 125 1461 MXI2XL $T=324800 470380 0 0 $X=324200 $Y=470020
X758 1238 1177 15 14 126 1463 MXI2XL $T=332920 418180 1 0 $X=332320 $Y=412360
X759 257 1180 15 14 798 254 MXI2XL $T=333500 522580 1 0 $X=332900 $Y=516760
X760 1492 1183 15 14 125 1518 MXI2XL $T=353220 459940 1 0 $X=352620 $Y=454120
X761 1519 1188 15 14 126 1520 MXI2XL $T=353800 397300 1 0 $X=353200 $Y=391480
X762 290 1190 15 14 125 280 MXI2XL $T=364240 459940 0 180 $X=359000 $Y=454120
X763 283 1191 15 14 125 1521 MXI2XL $T=369460 491260 0 180 $X=364220 $Y=485440
X764 1373 1192 15 14 126 1372 MXI2XL $T=371200 386860 0 0 $X=370600 $Y=386500
X765 289 1197 15 14 126 294 MXI2XL $T=386280 418180 0 0 $X=385680 $Y=417820
X766 1468 1201 15 14 798 311 MXI2XL $T=401360 522580 1 180 $X=396120 $Y=522220
X767 1398 1210 15 14 125 396 MXI2XL $T=473860 459940 0 180 $X=468620 $Y=454120
X768 176 1212 15 14 126 399 MXI2XL $T=481980 386860 1 180 $X=476740 $Y=386500
X769 1406 1253 15 14 797 1409 MXI2XL $T=485460 522580 0 0 $X=484860 $Y=522220
X770 1522 1214 15 14 125 1523 MXI2XL $T=490680 480820 1 180 $X=485440 $Y=480460
X771 1524 1215 15 14 126 1525 MXI2XL $T=497060 418180 1 180 $X=491820 $Y=417820
X772 1283 1220 15 14 125 1526 MXI2XL $T=498800 480820 0 180 $X=493560 $Y=475000
X773 1527 1222 15 14 125 401 MXI2XL $T=501700 449500 0 180 $X=496460 $Y=443680
X774 1285 1217 15 14 126 1482 MXI2XL $T=498220 407740 0 0 $X=497620 $Y=407380
X775 411 1219 15 14 798 409 MXI2XL $T=503440 522580 0 0 $X=502840 $Y=522220
X776 1485 1227 15 14 125 1261 MXI2XL $T=524900 491260 0 180 $X=519660 $Y=485440
X777 197 1234 15 14 126 1259 MXI2XL $T=530120 397300 0 180 $X=524880 $Y=391480
X778 1528 1529 15 14 1361 1521 AND3X1 $T=347420 491260 1 0 $X=346820 $Y=485440
X779 1530 1531 15 14 1363 294 AND3X1 $T=368300 418180 0 0 $X=367700 $Y=417820
X780 1468 797 15 14 1146 326 AND3X1 $T=403100 522580 0 0 $X=402500 $Y=522220
X781 1342 15 14 622 1341 1171 623 714 AOI221XL $T=318420 522580 1 180 $X=312020 $Y=522220
X782 253 15 14 1344 723 1532 629 125 AOI221XL $T=321320 470380 1 0 $X=320720 $Y=464560
X783 1238 15 14 1345 1174 1533 634 126 AOI221XL $T=332340 418180 0 180 $X=325940 $Y=412360
X784 723 15 14 639 1493 252 1352 1465 AOI221XL $T=331180 449500 0 0 $X=330580 $Y=449140
X785 723 15 14 701 283 1534 1367 125 AOI221XL $T=369460 491260 1 0 $X=368860 $Y=485440
X786 1174 15 14 694 289 1535 1369 126 AOI221XL $T=379900 418180 0 0 $X=379300 $Y=417820
X787 1261 15 14 1425 731 1536 818 129 AOI221XL $T=524900 480820 0 0 $X=524300 $Y=480460
X788 1259 15 14 1422 158 1537 199 135 AOI221XL $T=525480 397300 0 0 $X=524880 $Y=396940
X789 1286 302 15 14 303 1538 129 697 BMXIX2 $T=383960 491260 1 0 $X=383360 $Y=485440
X790 1288 304 15 14 305 1539 135 708 BMXIX2 $T=395560 428620 1 0 $X=394960 $Y=422800
X791 1277 347 15 14 346 1508 129 715 BMXIX2 $T=424560 480820 1 180 $X=408880 $Y=480460
X792 1501 347 15 14 346 1269 129 729 BMXIX2 $T=414120 480820 1 0 $X=413520 $Y=475000
X793 1281 355 15 14 354 1504 135 724 BMXIX2 $T=433260 418180 1 180 $X=417580 $Y=417820
X794 1506 355 15 14 354 1273 135 732 BMXIX2 $T=425140 418180 1 0 $X=424540 $Y=412360
X795 1297 388 15 14 389 1540 125 740 BMXIX2 $T=465160 501700 0 180 $X=449480 $Y=495880
X796 1251 387 15 14 386 1248 563 453 BMXIX2 $T=465740 533020 0 180 $X=450060 $Y=527200
X797 1294 394 15 14 395 1541 126 751 BMXIX2 $T=468060 407740 0 0 $X=467460 $Y=407380
X798 1542 437 15 14 34 491 ADDHX1 $T=52780 386860 0 0 $X=52180 $Y=386500
X799 1543 33 15 14 32 493 ADDHX1 $T=54520 376420 0 0 $X=53920 $Y=376060
X800 1544 492 15 14 469 495 ADDHX1 $T=62640 439060 0 0 $X=62040 $Y=438700
X801 1545 490 15 14 475 510 ADDHX1 $T=69020 418180 0 0 $X=68420 $Y=417820
X802 1546 494 15 14 484 515 ADDHX1 $T=93960 449500 0 180 $X=84080 $Y=443680
X803 1547 514 15 14 530 505 ADDHX1 $T=100920 407740 1 180 $X=91040 $Y=407380
X804 1548 509 15 14 499 539 ADDHX1 $T=96860 439060 1 0 $X=96260 $Y=433240
X805 1549 538 15 14 540 1035 ADDHX1 $T=152540 428620 1 0 $X=151940 $Y=422800
X806 1310 75 15 14 1043 1550 ADDHX1 $T=171680 386860 1 180 $X=161800 $Y=386500
X807 1551 1044 15 14 75 1552 ADDHX1 $T=188500 397300 0 180 $X=178620 $Y=391480
X808 1319 1106 15 14 1051 1553 ADDHX1 $T=223880 470380 0 0 $X=223280 $Y=470020
X809 1554 1052 15 14 1106 1555 ADDHX1 $T=224460 449500 1 0 $X=223860 $Y=443680
X810 1326 1138 15 14 1101 1556 ADDHX1 $T=252880 470380 1 0 $X=252280 $Y=464560
X811 1557 1102 15 14 1138 1558 ADDHX1 $T=288260 459940 1 0 $X=287660 $Y=454120
X812 1333 1095 15 14 1133 1559 ADDHX1 $T=289420 418180 0 0 $X=288820 $Y=417820
X813 1560 1134 15 14 1095 1561 ADDHX1 $T=301020 397300 0 180 $X=291140 $Y=391480
X814 1265 688 15 14 555 284 ADDHX1 $T=374680 533020 1 180 $X=364800 $Y=532660
X815 1496 706 15 14 722 302 ADDHX1 $T=392660 480820 0 0 $X=392060 $Y=480460
X816 316 1144 15 14 723 312 ADDHX1 $T=407740 491260 1 180 $X=397860 $Y=490900
X817 1498 718 15 14 1237 304 ADDHX1 $T=403680 418180 0 0 $X=403080 $Y=417820
X818 1562 1148 15 14 722 342 ADDHX1 $T=406000 491260 1 0 $X=405400 $Y=485440
X819 1301 721 15 14 1174 328 ADDHX1 $T=419920 428620 0 180 $X=410040 $Y=422800
X820 1563 754 15 14 1237 336 ADDHX1 $T=423980 418180 0 180 $X=414100 $Y=412360
X821 1303 1150 15 14 564 348 ADDHX1 $T=421080 533020 0 0 $X=420480 $Y=532660
X822 1305 1154 15 14 731 372 ADDHX1 $T=441380 491260 0 0 $X=440780 $Y=490900
X823 1307 742 15 14 158 364 ADDHX1 $T=453560 439060 0 180 $X=443680 $Y=433240
X824 1511 749 15 14 730 388 ADDHX1 $T=452400 480820 0 0 $X=451800 $Y=480460
X825 1513 756 15 14 1216 394 ADDHX1 $T=452980 407740 0 0 $X=452380 $Y=407380
X826 75 15 14 1030 237 1309 AO21X1 $T=170520 397300 1 0 $X=169920 $Y=391480
X827 1031 15 14 1044 75 1432 AO21X1 $T=201260 397300 0 0 $X=200660 $Y=396940
X828 1106 15 14 1026 241 1318 AO21X1 $T=215180 470380 0 0 $X=214580 $Y=470020
X829 1027 15 14 1052 1106 1437 AO21X1 $T=227940 459940 1 0 $X=227340 $Y=454120
X830 1138 15 14 1075 247 1325 AO21X1 $T=261000 480820 1 0 $X=260400 $Y=475000
X831 1076 15 14 1102 1138 1449 AO21X1 $T=275500 470380 1 0 $X=274900 $Y=464560
X832 1095 15 14 1129 249 1332 AO21X1 $T=291740 418180 1 0 $X=291140 $Y=412360
X833 1130 15 14 1134 1095 1453 AO21X1 $T=294640 407740 0 0 $X=294040 $Y=407380
X834 619 15 14 641 714 1460 AO21X1 $T=307980 512140 0 0 $X=307380 $Y=511780
X835 125 15 14 1564 1532 1172 AO21X1 $T=323060 470380 1 180 $X=317240 $Y=470020
X836 126 15 14 1565 1533 1176 AO21X1 $T=328280 407740 1 180 $X=322460 $Y=407380
X837 722 15 14 1343 252 258 AO21X1 $T=330600 470380 0 0 $X=330000 $Y=470020
X838 723 15 14 1343 1461 1566 AO21X1 $T=331180 470380 1 0 $X=330580 $Y=464560
X839 1529 15 14 1566 129 1567 AO21X1 $T=332920 480820 0 0 $X=332320 $Y=480460
X840 1174 15 14 1349 1463 1568 AO21X1 $T=342780 418180 0 180 $X=336960 $Y=412360
X841 1357 15 14 1569 129 1570 AO21X1 $T=337560 449500 0 0 $X=336960 $Y=449140
X842 657 15 14 723 1566 274 AO21X1 $T=338140 480820 0 0 $X=337540 $Y=480460
X843 657 15 14 722 258 1240 AO21X1 $T=339300 470380 0 0 $X=338700 $Y=470020
X844 654 15 14 723 1518 1569 AO21X1 $T=341620 449500 1 0 $X=341020 $Y=443680
X845 1358 15 14 1571 135 1572 AO21X1 $T=343360 397300 1 0 $X=342760 $Y=391480
X846 1531 15 14 1568 135 1573 AO21X1 $T=352640 418180 0 180 $X=346820 $Y=412360
X847 646 15 14 1174 1520 1571 AO21X1 $T=353800 397300 0 180 $X=347980 $Y=391480
X848 675 15 14 1237 262 1244 AO21X1 $T=352640 407740 0 0 $X=352040 $Y=407380
X849 675 15 14 1174 1568 276 AO21X1 $T=353800 418180 1 0 $X=353200 $Y=412360
X850 125 15 14 1574 1534 1193 AO21X1 $T=359600 491260 1 0 $X=359000 $Y=485440
X851 723 15 14 1366 1521 292 AO21X1 $T=366560 470380 0 0 $X=365960 $Y=470020
X852 722 15 14 1366 282 1575 AO21X1 $T=370620 480820 1 0 $X=370020 $Y=475000
X853 1237 15 14 296 288 1576 AO21X1 $T=378160 407740 0 0 $X=377560 $Y=407380
X854 301 15 14 1575 125 1577 AO21X1 $T=385120 480820 0 180 $X=379300 $Y=475000
X855 703 15 14 723 292 298 AO21X1 $T=384540 470380 0 0 $X=383940 $Y=470020
X856 703 15 14 722 1575 1287 AO21X1 $T=386280 480820 1 0 $X=385680 $Y=475000
X857 1141 15 14 695 714 1469 AO21X1 $T=386280 522580 1 0 $X=385680 $Y=516760
X858 126 15 14 1578 1535 1194 AO21X1 $T=386860 428620 1 0 $X=386260 $Y=422800
X859 709 15 14 1237 1576 1289 AO21X1 $T=395560 407740 1 180 $X=389740 $Y=407380
X860 722 15 14 1378 1466 314 AO21X1 $T=394980 459940 0 0 $X=394380 $Y=459580
X861 723 15 14 1378 300 1579 AO21X1 $T=394980 470380 0 0 $X=394380 $Y=470020
X862 309 15 14 1576 126 1580 AO21X1 $T=395560 407740 0 0 $X=394960 $Y=407380
X863 722 15 14 1379 1287 1581 AO21X1 $T=400780 480820 1 0 $X=400180 $Y=475000
X864 723 15 14 1379 298 1291 AO21X1 $T=402520 470380 1 0 $X=401920 $Y=464560
X865 1237 15 14 1381 1470 1271 AO21X1 $T=404260 397300 0 0 $X=403660 $Y=396940
X866 1174 15 14 1381 308 1582 AO21X1 $T=404260 407740 1 0 $X=403660 $Y=401920
X867 1237 15 14 345 1289 334 AO21X1 $T=420500 407740 1 180 $X=414680 $Y=407380
X868 1151 15 14 726 1251 1250 AO21X1 $T=423400 522580 0 0 $X=422800 $Y=522220
X869 731 15 14 1392 390 368 AO21X1 $T=451820 470380 1 180 $X=446000 $Y=470020
X870 730 15 14 1392 1299 366 AO21X1 $T=452400 480820 1 180 $X=446580 $Y=480460
X871 1216 15 14 1395 1296 378 AO21X1 $T=460520 418180 1 180 $X=454700 $Y=417820
X872 730 15 14 1399 1477 1275 AO21X1 $T=468060 480820 1 0 $X=467460 $Y=475000
X873 761 15 14 730 1583 1299 AO21X1 $T=477340 480820 1 180 $X=471520 $Y=480460
X874 1216 15 14 1400 1481 1279 AO21X1 $T=472700 418180 0 0 $X=472100 $Y=417820
X875 759 15 14 1216 1584 1296 AO21X1 $T=474440 428620 1 0 $X=473840 $Y=422800
X876 765 15 14 768 728 1479 AO21X1 $T=477340 522580 1 0 $X=476740 $Y=516760
X877 1298 15 14 1583 129 1585 AO21X1 $T=483720 480820 0 180 $X=477900 $Y=475000
X878 1295 15 14 1584 135 1586 AO21X1 $T=479660 418180 0 0 $X=479060 $Y=417820
X879 764 15 14 767 728 1480 AO21X1 $T=482560 522580 1 0 $X=481960 $Y=516760
X880 1216 15 14 404 1482 1584 AO21X1 $T=488360 407740 1 180 $X=482540 $Y=407380
X881 730 15 14 402 1526 1583 AO21X1 $T=492420 480820 0 180 $X=486600 $Y=475000
X882 186 15 14 1216 406 413 AO21X1 $T=499960 376420 0 0 $X=499360 $Y=376060
X883 773 15 14 731 1527 1587 AO21X1 $T=500540 439060 0 0 $X=499940 $Y=438700
X884 773 15 14 730 400 423 AO21X1 $T=501700 449500 1 0 $X=501100 $Y=443680
X885 795 15 14 806 728 1483 AO21X1 $T=508080 522580 1 0 $X=507480 $Y=516760
X886 193 15 14 187 126 1588 AO21X1 $T=513880 376420 1 180 $X=508060 $Y=376060
X887 189 15 14 1216 429 1255 AO21X1 $T=515040 397300 1 180 $X=509220 $Y=396940
X888 435 15 14 1589 126 1590 AO21X1 $T=515620 407740 0 180 $X=509800 $Y=401920
X889 1414 15 14 1587 125 1591 AO21X1 $T=510980 439060 0 0 $X=510380 $Y=438700
X890 794 15 14 805 728 1484 AO21X1 $T=510980 512140 0 0 $X=510380 $Y=511780
X891 189 15 14 158 1589 1592 AO21X1 $T=511560 397300 1 0 $X=510960 $Y=391480
X892 1421 15 14 1593 129 1594 AO21X1 $T=517360 470380 1 180 $X=511540 $Y=470020
X893 799 15 14 730 1593 1595 AO21X1 $T=513300 470380 1 0 $X=512700 $Y=464560
X894 799 15 14 731 431 1596 AO21X1 $T=513880 480820 0 0 $X=513280 $Y=480460
X895 158 15 14 196 197 1589 AO21X1 $T=518520 397300 1 0 $X=517920 $Y=391480
X896 731 15 14 1424 1485 431 AO21X1 $T=524900 480820 1 180 $X=519080 $Y=480460
X897 129 15 14 1597 1536 1233 AO21X1 $T=530700 480820 0 0 $X=530100 $Y=480460
X898 135 15 14 1598 1537 1228 AO21X1 $T=531280 397300 0 0 $X=530680 $Y=396940
X899 72 1550 15 14 1426 XNOR2X1 $T=161240 386860 1 0 $X=160640 $Y=381040
X900 74 1552 15 14 1487 XNOR2X1 $T=179220 386860 0 0 $X=178620 $Y=386500
X901 92 84 15 14 1034 XNOR2X1 $T=217500 376420 0 0 $X=216900 $Y=376060
X902 1045 1555 15 14 1488 XNOR2X1 $T=231420 449500 1 180 $X=224440 $Y=449140
X903 1046 1553 15 14 1434 XNOR2X1 $T=239540 470380 1 180 $X=232560 $Y=470020
X904 1135 1556 15 14 1443 XNOR2X1 $T=274340 470380 0 180 $X=267360 $Y=464560
X905 1124 1561 15 14 1489 XNOR2X1 $T=288260 386860 0 0 $X=287660 $Y=386500
X906 1136 1558 15 14 1490 XNOR2X1 $T=291740 449500 0 0 $X=291140 $Y=449140
X907 1123 1559 15 14 1456 XNOR2X1 $T=299860 418180 0 0 $X=299260 $Y=417820
X908 286 680 15 14 555 XNOR2X1 $T=372940 522580 1 180 $X=365960 $Y=522220
X909 669 734 15 14 682 XNOR2X1 $T=369460 470380 1 0 $X=368860 $Y=464560
X910 684 692 15 14 736 XNOR2X1 $T=392080 386860 1 180 $X=385100 $Y=386500
X911 340 564 15 14 555 XNOR2X1 $T=416440 533020 1 180 $X=409460 $Y=532660
X912 346 730 15 14 723 XNOR2X1 $T=424560 491260 0 180 $X=417580 $Y=485440
X913 354 1216 15 14 1174 XNOR2X1 $T=428620 428620 1 0 $X=428020 $Y=422800
X914 350 560 15 14 731 XNOR2X1 $T=437900 501700 1 0 $X=437300 $Y=495880
X915 561 737 15 14 158 XNOR2X1 $T=452980 428620 1 180 $X=446000 $Y=428260
X916 386 455 15 14 728 XNOR2X1 $T=459360 522580 1 180 $X=452380 $Y=522220
X917 748 755 15 14 752 XNOR2X1 $T=456460 397300 1 0 $X=455860 $Y=391480
X918 758 744 15 14 746 XNOR2X1 $T=457620 459940 0 0 $X=457020 $Y=459580
X919 125 15 14 260 259 1567 1181 OAI31XL $T=339880 480820 0 180 $X=334640 $Y=475000
X920 125 15 14 1465 1493 1570 1178 OAI31XL $T=342780 459940 0 180 $X=337540 $Y=454120
X921 648 15 14 666 554 555 254 OAI31XL $T=344520 522580 0 180 $X=339280 $Y=516760
X922 126 15 14 270 263 1573 1185 OAI31XL $T=346260 407740 0 0 $X=345660 $Y=407380
X923 126 15 14 268 273 1572 1175 OAI31XL $T=351480 397300 1 180 $X=346240 $Y=396940
X924 129 15 14 1466 293 1577 1195 OAI31XL $T=379900 470380 0 0 $X=379300 $Y=470020
X925 135 15 14 1470 1494 1580 1199 OAI31XL $T=400780 407740 0 0 $X=400180 $Y=407380
X926 1471 15 14 323 1599 1600 1202 OAI31XL $T=408900 480820 1 0 $X=408300 $Y=475000
X927 1268 15 14 314 324 125 1600 OAI31XL $T=415860 470380 0 180 $X=410620 $Y=464560
X928 1272 15 14 1271 352 126 1601 OAI31XL $T=431520 407740 1 0 $X=430920 $Y=401920
X929 1472 15 14 333 1602 1601 1206 OAI31XL $T=434420 407740 0 0 $X=433820 $Y=407380
X930 1276 15 14 1275 358 129 1603 OAI31XL $T=434420 480820 1 0 $X=433820 $Y=475000
X931 1473 15 14 371 1604 1603 1204 OAI31XL $T=440220 491260 0 180 $X=434980 $Y=485440
X932 1474 15 14 383 1605 1606 1205 OAI31XL $T=443700 428620 0 180 $X=438460 $Y=422800
X933 1280 15 14 1279 362 135 1606 OAI31XL $T=444280 418180 1 180 $X=439040 $Y=417820
X934 125 15 14 1477 1517 1585 1211 OAI31XL $T=477340 480820 0 0 $X=476740 $Y=480460
X935 126 15 14 1481 1516 1586 1209 OAI31XL $T=480820 418180 1 0 $X=480220 $Y=412360
X936 135 15 14 417 414 1588 1231 OAI31XL $T=507500 386860 1 0 $X=506900 $Y=381040
X937 125 15 14 420 432 1594 1225 OAI31XL $T=511560 491260 1 0 $X=510960 $Y=485440
X938 129 15 14 427 424 1591 1229 OAI31XL $T=512140 449500 1 0 $X=511540 $Y=443680
X939 135 15 14 425 430 1590 1226 OAI31XL $T=515620 407740 1 0 $X=515020 $Y=401920
X940 1529 1361 15 14 274 129 1360 AOI31XL $T=340460 491260 1 0 $X=339860 $Y=485440
X941 554 648 15 14 666 714 256 AOI31XL $T=345100 512140 1 180 $X=339860 $Y=511780
X942 1531 1363 15 14 276 135 1365 AOI31XL $T=361340 418180 0 0 $X=360740 $Y=417820
X943 461 455 15 14 562 728 1416 AOI31XL $T=472120 522580 1 0 $X=471520 $Y=516760
X944 419 407 15 14 1596 125 1411 AOI31XL $T=513300 480820 1 180 $X=508060 $Y=480460
X945 435 434 15 14 1592 126 1413 AOI31XL $T=517940 407740 1 180 $X=512700 $Y=407380
X946 1315 1312 15 14 1157 1429 1313 AOI211XL $T=204160 386860 0 180 $X=199500 $Y=381040
X947 1324 1321 15 14 1160 1441 1322 AOI211XL $T=245920 449500 0 0 $X=245320 $Y=449140
X948 1328 1329 15 14 1167 1448 1330 AOI211XL $T=280140 459940 0 0 $X=279540 $Y=459580
X949 1340 1337 15 14 1164 1455 1338 AOI211XL $T=302180 397300 0 0 $X=301580 $Y=396940
X950 704 722 15 14 1538 1466 299 AOI211XL $T=392080 470380 0 180 $X=387420 $Y=464560
X951 710 1237 15 14 1539 1470 1497 AOI211XL $T=399620 397300 0 0 $X=399020 $Y=396940
X952 1385 1599 15 14 1500 1471 1579 AOI211XL $T=412960 470380 1 180 $X=408300 $Y=470020
X953 721 1237 15 14 1302 1271 1502 AOI211XL $T=415860 407740 1 0 $X=415260 $Y=401920
X954 1389 1602 15 14 1505 1472 1582 AOI211XL $T=433260 407740 1 180 $X=428600 $Y=407380
X955 1386 1605 15 14 1503 1474 1476 AOI211XL $T=435000 428620 1 0 $X=434400 $Y=422800
X956 1387 1604 15 14 1507 1473 1475 AOI211XL $T=435000 480820 0 0 $X=434400 $Y=480460
X957 1154 730 15 14 1306 1275 369 AOI211XL $T=443120 480820 1 0 $X=442520 $Y=475000
X958 742 1216 15 14 1308 1279 375 AOI211XL $T=448340 418180 0 0 $X=447740 $Y=417820
X959 762 730 15 14 1540 1477 391 AOI211XL $T=460520 491260 1 0 $X=459920 $Y=485440
X960 760 1216 15 14 1541 1481 1514 AOI211XL $T=475600 418180 0 180 $X=470940 $Y=412360
X961 322 15 14 317 1581 318 1290 125 AOI32XL $T=401940 480820 0 0 $X=401340 $Y=480460
X962 628 15 14 723 1564 1461 ACHCONX2 $T=305660 459940 0 0 $X=305080 $Y=459580
X963 633 15 14 1174 1565 1463 ACHCONX2 $T=311460 407740 1 0 $X=310880 $Y=401920
X964 631 15 14 1174 1464 1571 ACHCONX2 $T=313200 386860 0 0 $X=312620 $Y=386500
X965 638 15 14 723 1462 1569 ACHCONX2 $T=318420 439060 0 0 $X=317840 $Y=438700
X966 661 15 14 722 1528 275 ACHCONX2 $T=324800 491260 0 0 $X=324220 $Y=490900
X967 674 15 14 716 1520 1372 ACHCONX2 $T=342200 386860 0 0 $X=341620 $Y=386500
X968 678 15 14 1237 1530 277 ACHCONX2 $T=344520 428620 1 0 $X=343940 $Y=422800
X969 664 15 14 722 1518 281 ACHCONX2 $T=346260 449500 0 0 $X=345680 $Y=449140
X970 716 15 14 673 1519 1373 ACHCONX2 $T=346840 386860 1 0 $X=346260 $Y=381040
X971 663 15 14 722 1492 291 ACHCONX2 $T=346840 449500 1 0 $X=346260 $Y=443680
X972 700 15 14 723 1574 1521 ACHCONX2 $T=375840 480820 1 180 $X=346260 $Y=480460
X973 693 15 14 1174 1578 294 ACHCONX2 $T=407160 418180 0 180 $X=377580 $Y=412360
X974 743 15 14 723 1267 325 ACHCONX2 $T=436740 449500 1 180 $X=407160 $Y=449140
X975 733 15 14 731 1274 359 ACHCONX2 $T=417020 470380 1 0 $X=416440 $Y=464560
X976 716 15 14 158 1278 363 ACHCONX2 $T=417600 428620 0 0 $X=417020 $Y=428260
X977 160 15 14 1174 1270 353 ACHCONX2 $T=448920 397300 1 180 $X=419340 $Y=396940
X978 175 15 14 162 406 398 ACHCONX2 $T=468060 376420 0 0 $X=467480 $Y=376060
X979 458 15 14 397 400 731 ACHCONX2 $T=468060 449500 1 0 $X=467480 $Y=443680
X980 458 15 14 730 1527 1398 ACHCONX2 $T=468060 449500 0 0 $X=467480 $Y=449140
X981 770 15 14 730 1523 1526 ACHCONX2 $T=468060 470380 0 0 $X=467480 $Y=470020
X982 781 15 14 1216 1525 1482 ACHCONX2 $T=471540 407740 1 0 $X=470960 $Y=401920
X983 771 15 14 730 1522 1283 ACHCONX2 $T=476180 491260 1 0 $X=475600 $Y=485440
X984 782 15 14 1216 1524 1285 ACHCONX2 $T=485460 418180 1 0 $X=484880 $Y=412360
X985 791 15 14 731 1282 1596 ACHCONX2 $T=488940 459940 0 0 $X=488360 $Y=459580
X986 789 15 14 158 1284 1592 ACHCONX2 $T=498800 418180 0 0 $X=498220 $Y=417820
X987 802 15 14 731 1486 1587 ACHCONX2 $T=533600 439060 0 180 $X=504020 $Y=433240
X988 192 15 14 158 1598 197 ACHCONX2 $T=512140 386860 0 0 $X=511560 $Y=386500
X989 194 15 14 158 203 187 ACHCONX2 $T=513880 376420 0 0 $X=513300 $Y=376060
X990 817 15 14 731 1597 1485 ACHCONX2 $T=516780 480820 1 0 $X=516200 $Y=475000
X991 1240 15 14 261 1243 129 1359 AND4XL $T=349740 480820 0 180 $X=343920 $Y=475000
X992 1244 15 14 271 1247 135 1364 AND4XL $T=361340 407740 0 0 $X=360740 $Y=407380
X993 1595 15 14 1421 416 125 1410 AND4XL $T=510980 470380 1 180 $X=505160 $Y=470020
X994 1255 15 14 426 1257 126 1412 AND4XL $T=511560 407740 1 180 $X=505740 $Y=407380
X995 1607 15 14 573 28 1608 470 ADDFXL $T=54520 407740 1 180 $X=38840 $Y=407380
X996 1609 15 14 568 576 1610 827 ADDFXL $T=55100 480820 1 180 $X=39420 $Y=480460
X997 1608 15 14 565 32 1611 473 ADDFXL $T=41760 397300 0 0 $X=41160 $Y=396940
X998 1612 15 14 571 570 1613 831 ADDFXL $T=57420 501700 1 180 $X=41740 $Y=501340
X999 1613 15 14 575 574 1614 843 ADDFXL $T=42920 428620 1 0 $X=42320 $Y=422800
X1000 1610 15 14 570 578 1615 823 ADDFXL $T=58000 449500 1 180 $X=42320 $Y=449140
X1001 1614 15 14 577 566 31 477 ADDFXL $T=43500 407740 1 0 $X=42900 $Y=401920
X1002 1616 15 14 569 578 1607 822 ADDFXL $T=58580 459940 0 180 $X=42900 $Y=454120
X1003 1617 15 14 567 576 1616 826 ADDFXL $T=58580 480820 0 180 $X=42900 $Y=475000
X1004 1618 15 14 572 570 1619 830 ADDFXL $T=58580 501700 0 180 $X=42900 $Y=495880
X1005 1620 15 14 578 566 1621 476 ADDFXL $T=44080 418180 1 0 $X=43480 $Y=412360
X1006 1622 15 14 579 568 1612 835 ADDFXL $T=59160 543460 0 180 $X=43480 $Y=537640
X1007 1619 15 14 576 574 1620 842 ADDFXL $T=44660 428620 0 0 $X=44060 $Y=428260
X1008 1623 15 14 582 572 1609 839 ADDFXL $T=59740 522580 1 180 $X=44060 $Y=522220
X1009 1624 15 14 581 572 1617 838 ADDFXL $T=59740 533020 1 180 $X=44060 $Y=532660
X1010 1625 15 14 580 568 1618 834 ADDFXL $T=60900 533020 0 180 $X=45220 $Y=527200
X1011 1621 15 14 28 34 1543 41 ADDFXL $T=51040 386860 1 0 $X=50440 $Y=381040
X1012 1626 15 14 566 32 1542 474 ADDFXL $T=52200 397300 1 0 $X=51600 $Y=391480
X1013 1615 15 14 574 28 1626 471 ADDFXL $T=54520 407740 0 0 $X=53920 $Y=407380
X1014 1627 15 14 828 469 1628 479 ADDFXL $T=55100 480820 0 0 $X=54500 $Y=480460
X1015 1629 15 14 829 469 1630 480 ADDFXL $T=70180 491260 0 180 $X=54500 $Y=485440
X1016 1631 15 14 821 36 1544 488 ADDFXL $T=71920 459940 1 180 $X=56240 $Y=459580
X1017 1632 15 14 833 821 1629 486 ADDFXL $T=75980 501700 0 180 $X=60300 $Y=495880
X1018 1633 15 14 832 821 1627 485 ADDFXL $T=75980 501700 1 180 $X=60300 $Y=501340
X1019 1634 15 14 836 841 1635 501 ADDFXL $T=76560 470380 1 180 $X=60880 $Y=470020
X1020 1630 15 14 841 472 1545 498 ADDFXL $T=62640 439060 1 0 $X=62040 $Y=433240
X1021 1636 15 14 820 36 1637 489 ADDFXL $T=64960 449500 1 0 $X=64360 $Y=443680
X1022 1628 15 14 840 472 1638 497 ADDFXL $T=65540 428620 0 0 $X=64940 $Y=428260
X1023 1635 15 14 824 475 1636 483 ADDFXL $T=65540 470380 1 0 $X=64940 $Y=464560
X1024 1639 15 14 585 580 1624 850 ADDFXL $T=65540 533020 0 0 $X=64940 $Y=532660
X1025 1640 15 14 583 582 1622 847 ADDFXL $T=65540 543460 0 0 $X=64940 $Y=543100
X1026 1641 15 14 584 582 1625 846 ADDFXL $T=66120 543460 1 0 $X=65520 $Y=537640
X1027 1642 15 14 586 580 1623 851 ADDFXL $T=66700 533020 1 0 $X=66100 $Y=527200
X1028 1643 15 14 844 825 1633 854 ADDFXL $T=82940 512140 0 180 $X=67260 $Y=506320
X1029 1644 15 14 837 841 1645 500 ADDFXL $T=70180 480820 0 0 $X=69580 $Y=480460
X1030 1646 15 14 848 829 1634 862 ADDFXL $T=70180 491260 1 0 $X=69580 $Y=485440
X1031 1645 15 14 825 475 1631 482 ADDFXL $T=71920 459940 0 0 $X=71320 $Y=459580
X1032 1647 15 14 849 829 1644 861 ADDFXL $T=75980 501700 1 0 $X=75380 $Y=495880
X1033 1648 15 14 845 825 1632 855 ADDFXL $T=75980 501700 0 0 $X=75380 $Y=501340
X1034 1649 15 14 853 487 1546 503 ADDFXL $T=100340 449500 1 180 $X=84660 $Y=449140
X1035 1650 15 14 587 586 1640 874 ADDFXL $T=86420 543460 0 0 $X=85820 $Y=543100
X1036 1651 15 14 852 487 1652 504 ADDFXL $T=102080 459940 1 180 $X=86400 $Y=459580
X1037 1653 15 14 867 481 1651 513 ADDFXL $T=102080 470380 0 180 $X=86400 $Y=464560
X1038 1654 15 14 588 586 1641 873 ADDFXL $T=87000 533020 0 0 $X=86400 $Y=532660
X1039 1655 15 14 589 584 1639 877 ADDFXL $T=87000 543460 1 0 $X=86400 $Y=537640
X1040 1656 15 14 590 584 1642 878 ADDFXL $T=87580 533020 1 0 $X=86980 $Y=527200
X1041 1657 15 14 875 833 1646 866 ADDFXL $T=103820 512140 0 180 $X=88140 $Y=506320
X1042 1658 15 14 871 837 1643 869 ADDFXL $T=88740 512140 0 0 $X=88140 $Y=511780
X1043 1659 15 14 48 506 1660 47 ADDFXL $T=106140 386860 0 180 $X=90460 $Y=381040
X1044 1661 15 14 860 496 1548 527 ADDFXL $T=106140 439060 1 180 $X=90460 $Y=438700
X1045 1662 15 14 868 481 1649 512 ADDFXL $T=106140 459940 0 180 $X=90460 $Y=454120
X1046 1663 15 14 876 833 1647 865 ADDFXL $T=106140 501700 0 180 $X=90460 $Y=495880
X1047 1664 15 14 872 837 1648 870 ADDFXL $T=91060 501700 0 0 $X=90460 $Y=501340
X1048 1665 15 14 927 506 1666 50 ADDFXL $T=123540 397300 0 180 $X=107860 $Y=391480
X1049 1667 15 14 892 502 1547 507 ADDFXL $T=123540 407740 1 180 $X=107860 $Y=407380
X1050 1668 15 14 891 502 1669 508 ADDFXL $T=123540 418180 0 180 $X=107860 $Y=412360
X1051 1670 15 14 859 496 1671 526 ADDFXL $T=108460 449500 1 0 $X=107860 $Y=443680
X1052 1672 15 14 888 484 1673 524 ADDFXL $T=123540 459940 1 180 $X=107860 $Y=459580
X1053 1673 15 14 864 478 1661 518 ADDFXL $T=108460 470380 1 0 $X=107860 $Y=464560
X1054 1674 15 14 863 478 1670 517 ADDFXL $T=108460 470380 0 0 $X=107860 $Y=470020
X1055 1675 15 14 592 590 1654 885 ADDFXL $T=123540 533020 1 180 $X=107860 $Y=532660
X1056 63 15 14 57 519 1659 857 ADDFXL $T=125280 376420 1 180 $X=109600 $Y=376060
X1057 1676 15 14 594 588 1656 882 ADDFXL $T=110200 533020 1 0 $X=109600 $Y=527200
X1058 1677 15 14 593 588 1655 881 ADDFXL $T=110200 543460 1 0 $X=109600 $Y=537640
X1059 1678 15 14 880 845 1663 889 ADDFXL $T=110780 501700 0 0 $X=110180 $Y=501340
X1060 1679 15 14 879 845 1657 890 ADDFXL $T=111360 512140 1 0 $X=110760 $Y=506320
X1061 1680 15 14 591 590 1650 886 ADDFXL $T=126440 543460 1 180 $X=110760 $Y=543100
X1062 1681 15 14 887 484 1674 523 ADDFXL $T=127600 480820 0 180 $X=111920 $Y=475000
X1063 1682 15 14 911 511 1668 521 ADDFXL $T=129920 418180 1 180 $X=114240 $Y=417820
X1064 1683 15 14 915 868 1684 893 ADDFXL $T=131080 480820 1 180 $X=115400 $Y=480460
X1065 1685 15 14 923 533 1682 529 ADDFXL $T=131660 428620 0 180 $X=115980 $Y=422800
X1066 1686 15 14 883 849 1658 897 ADDFXL $T=117160 512140 0 0 $X=116560 $Y=511780
X1067 1687 15 14 884 849 1664 898 ADDFXL $T=117740 501700 1 0 $X=117140 $Y=495880
X1068 1688 15 14 930 519 1665 858 ADDFXL $T=133980 386860 1 180 $X=118300 $Y=386500
X1069 66 15 14 935 59 1688 49 ADDFXL $T=138620 386860 0 180 $X=122940 $Y=381040
X1070 1689 15 14 912 511 1667 520 ADDFXL $T=138620 407740 1 180 $X=122940 $Y=407380
X1071 1690 15 14 924 533 1689 528 ADDFXL $T=138620 418180 0 180 $X=122940 $Y=412360
X1072 1691 15 14 908 853 1672 532 ADDFXL $T=138620 459940 1 180 $X=122940 $Y=459580
X1073 1692 15 14 895 499 1653 535 ADDFXL $T=123540 470380 1 0 $X=122940 $Y=464560
X1074 1684 15 14 907 853 1681 531 ADDFXL $T=123540 470380 0 0 $X=122940 $Y=470020
X1075 1693 15 14 596 594 1675 901 ADDFXL $T=138620 533020 1 180 $X=122940 $Y=532660
X1076 1694 15 14 904 872 1678 909 ADDFXL $T=127020 501700 0 0 $X=126420 $Y=501340
X1077 1695 15 14 896 499 1662 534 ADDFXL $T=127600 459940 1 0 $X=127000 $Y=454120
X1078 1696 15 14 597 592 1677 905 ADDFXL $T=129340 543460 1 0 $X=128740 $Y=537640
X1079 1697 15 14 946 540 1685 537 ADDFXL $T=145000 418180 1 180 $X=129320 $Y=417820
X1080 1698 15 14 954 896 1683 913 ADDFXL $T=129920 480820 1 0 $X=129320 $Y=475000
X1081 1699 15 14 903 872 1679 910 ADDFXL $T=129920 512140 1 0 $X=129320 $Y=506320
X1082 1700 15 14 595 594 1680 902 ADDFXL $T=146740 543460 1 180 $X=131060 $Y=543100
X1083 1701 15 14 899 876 1686 921 ADDFXL $T=133400 522580 1 0 $X=132800 $Y=516760
X1084 1702 15 14 955 896 1703 914 ADDFXL $T=138620 459940 0 0 $X=138020 $Y=459580
X1085 1703 15 14 916 868 1691 894 ADDFXL $T=138620 470380 1 0 $X=138020 $Y=464560
X1086 1704 15 14 919 860 1692 542 ADDFXL $T=138620 470380 0 0 $X=138020 $Y=470020
X1087 1705 15 14 598 592 1676 906 ADDFXL $T=138620 533020 0 0 $X=138020 $Y=532660
X1088 1706 15 14 947 540 1690 536 ADDFXL $T=154280 418180 0 180 $X=138600 $Y=412360
X1089 1707 15 14 1031 947 1708 937 ADDFXL $T=155440 397300 0 180 $X=139760 $Y=391480
X1090 1709 15 14 938 884 1699 918 ADDFXL $T=155440 512140 1 180 $X=139760 $Y=511780
X1091 1710 15 14 999 912 1711 929 ADDFXL $T=156020 407740 1 180 $X=140340 $Y=407380
X1092 1712 15 14 998 912 1713 928 ADDFXL $T=156600 428620 1 180 $X=140920 $Y=428260
X1093 1714 15 14 900 876 1687 922 ADDFXL $T=141520 501700 1 0 $X=140920 $Y=495880
X1094 1715 15 14 920 860 1695 541 ADDFXL $T=157760 459940 0 180 $X=142080 $Y=454120
X1095 1716 15 14 939 884 1694 917 ADDFXL $T=158340 501700 1 180 $X=142660 $Y=501340
X1096 1717 15 14 601 596 1696 940 ADDFXL $T=144420 543460 1 0 $X=143820 $Y=537640
X1097 1718 15 14 994 924 1712 931 ADDFXL $T=160080 418180 1 180 $X=144400 $Y=417820
X1098 1708 15 14 995 924 1710 932 ADDFXL $T=149060 407740 1 0 $X=148460 $Y=401920
X1099 1719 15 14 943 880 1714 961 ADDFXL $T=150220 512140 1 0 $X=149620 $Y=506320
X1100 1720 15 14 974 920 1698 925 ADDFXL $T=165880 480820 0 180 $X=150200 $Y=475000
X1101 1721 15 14 942 880 1701 960 ADDFXL $T=150800 522580 1 0 $X=150200 $Y=516760
X1102 1722 15 14 599 598 1700 945 ADDFXL $T=150800 543460 0 0 $X=150200 $Y=543100
X1103 1723 15 14 602 596 1705 941 ADDFXL $T=153700 533020 0 0 $X=153100 $Y=532660
X1104 1724 15 14 1030 947 1718 936 ADDFXL $T=170520 397300 0 180 $X=154840 $Y=391480
X1105 1725 15 14 975 920 1702 926 ADDFXL $T=170520 459940 1 180 $X=154840 $Y=459580
X1106 1726 15 14 958 864 1704 953 ADDFXL $T=156020 470380 0 0 $X=155420 $Y=470020
X1107 1727 15 14 991 888 1728 980 ADDFXL $T=156600 470380 1 0 $X=156000 $Y=464560
X1108 1729 15 14 990 888 1726 981 ADDFXL $T=156600 480820 0 0 $X=156000 $Y=480460
X1109 1728 15 14 959 864 1715 952 ADDFXL $T=157760 459940 1 0 $X=157160 $Y=454120
X1110 1730 15 14 1044 1023 1707 934 ADDFXL $T=174580 397300 1 180 $X=158900 $Y=396940
X1111 1713 15 14 1002 892 1731 543 ADDFXL $T=159500 428620 0 0 $X=158900 $Y=428260
X1112 1732 15 14 966 900 1709 957 ADDFXL $T=159500 512140 0 0 $X=158900 $Y=511780
X1113 1733 15 14 600 598 1693 944 ADDFXL $T=159500 543460 1 0 $X=158900 $Y=537640
X1114 1711 15 14 1003 892 1734 544 ADDFXL $T=160080 418180 0 0 $X=159480 $Y=417820
X1115 1735 15 14 950 525 1736 545 ADDFXL $T=160660 439060 1 0 $X=160060 $Y=433240
X1116 1737 15 14 967 900 1716 956 ADDFXL $T=160660 501700 0 0 $X=160060 $Y=501340
X1117 1738 15 14 951 525 1549 546 ADDFXL $T=161820 428620 1 0 $X=161220 $Y=422800
X1118 1739 15 14 1043 1023 1724 933 ADDFXL $T=179220 407740 0 180 $X=163540 $Y=401920
X1119 1740 15 14 1010 959 1720 948 ADDFXL $T=180960 480820 0 180 $X=165280 $Y=475000
X1120 1741 15 14 971 904 1719 993 ADDFXL $T=165880 512140 1 0 $X=165280 $Y=506320
X1121 1742 15 14 970 904 1721 992 ADDFXL $T=165880 522580 1 0 $X=165280 $Y=516760
X1122 1743 15 14 603 600 1717 968 ADDFXL $T=165880 543460 0 0 $X=165280 $Y=543100
X1123 1744 15 14 963 908 1727 984 ADDFXL $T=173420 470380 1 0 $X=172820 $Y=464560
X1124 1745 15 14 978 516 1735 551 ADDFXL $T=174580 439060 0 0 $X=173980 $Y=438700
X1125 1746 15 14 606 602 1733 972 ADDFXL $T=174580 533020 0 0 $X=173980 $Y=532660
X1126 1747 15 14 604 600 1723 969 ADDFXL $T=174580 543460 1 0 $X=173980 $Y=537640
X1127 1748 15 14 1011 959 1725 949 ADDFXL $T=191400 459940 1 180 $X=175720 $Y=459580
X1128 1734 15 14 987 530 1749 548 ADDFXL $T=176900 418180 1 0 $X=176300 $Y=412360
X1129 1750 15 14 979 516 1738 552 ADDFXL $T=176900 428620 1 0 $X=176300 $Y=422800
X1130 1731 15 14 986 530 1751 547 ADDFXL $T=176900 428620 0 0 $X=176300 $Y=428260
X1131 1751 15 14 982 522 1745 549 ADDFXL $T=176900 439060 1 0 $X=176300 $Y=433240
X1132 1752 15 14 1019 943 1737 976 ADDFXL $T=178060 501700 0 0 $X=177460 $Y=501340
X1133 1753 15 14 1018 943 1732 977 ADDFXL $T=178060 512140 0 0 $X=177460 $Y=511780
X1134 236 15 14 1098 995 1754 81 ADDFXL $T=179220 407740 1 0 $X=178620 $Y=401920
X1135 1749 15 14 983 522 1750 550 ADDFXL $T=179220 418180 0 0 $X=178620 $Y=417820
X1136 1755 15 14 1007 916 1744 988 ADDFXL $T=179220 470380 0 0 $X=178620 $Y=470020
X1137 1756 15 14 1006 916 1757 989 ADDFXL $T=180380 491260 1 0 $X=179780 $Y=485440
X1138 238 15 14 75 995 1758 82 ADDFXL $T=180960 397300 0 0 $X=180360 $Y=396940
X1139 1757 15 14 962 908 1729 985 ADDFXL $T=180960 480820 1 0 $X=180360 $Y=475000
X1140 1759 15 14 1015 939 1741 965 ADDFXL $T=196040 512140 0 180 $X=180360 $Y=506320
X1141 1760 15 14 1014 939 1742 964 ADDFXL $T=196040 522580 0 180 $X=180360 $Y=516760
X1142 1761 15 14 605 602 1722 973 ADDFXL $T=180960 543460 0 0 $X=180360 $Y=543100
X1143 1758 15 14 1126 999 1762 87 ADDFXL $T=198360 407740 1 0 $X=197760 $Y=401920
X1144 1754 15 14 1125 999 1763 86 ADDFXL $T=198360 418180 1 0 $X=197760 $Y=412360
X1145 242 15 14 1114 1011 1764 996 ADDFXL $T=198360 459940 1 0 $X=197760 $Y=454120
X1146 1764 15 14 1102 975 1765 1000 ADDFXL $T=198360 459940 0 0 $X=197760 $Y=459580
X1147 1765 15 14 1076 955 1755 1004 ADDFXL $T=198360 470380 1 0 $X=197760 $Y=464560
X1148 240 15 14 1113 1011 1766 997 ADDFXL $T=198360 470380 0 0 $X=197760 $Y=470020
X1149 1766 15 14 1101 975 1767 1001 ADDFXL $T=198360 480820 1 0 $X=197760 $Y=475000
X1150 1767 15 14 1075 955 1756 1005 ADDFXL $T=198360 480820 0 0 $X=197760 $Y=480460
X1151 1768 15 14 608 606 1747 1021 ADDFXL $T=198360 543460 1 0 $X=197760 $Y=537640
X1152 1769 15 14 607 606 1743 1020 ADDFXL $T=198360 553900 1 0 $X=197760 $Y=548080
X1153 1770 15 14 1036 971 1753 1013 ADDFXL $T=198940 512140 0 0 $X=198340 $Y=511780
X1154 1771 15 14 610 604 1746 1016 ADDFXL $T=198940 533020 0 0 $X=198340 $Y=532660
X1155 1772 15 14 609 604 1761 1017 ADDFXL $T=198940 543460 0 0 $X=198340 $Y=543100
X1156 1773 15 14 1037 971 1752 1012 ADDFXL $T=200100 501700 0 0 $X=199500 $Y=501340
X1157 1774 15 14 1047 967 1760 1008 ADDFXL $T=200100 522580 1 0 $X=199500 $Y=516760
X1158 1775 15 14 1048 967 1759 1009 ADDFXL $T=201840 512140 1 0 $X=201240 $Y=506320
X1159 1776 15 14 1023 951 1706 1041 ADDFXL $T=213440 418180 1 0 $X=212840 $Y=412360
X1160 1777 15 14 1027 991 1748 1025 ADDFXL $T=228520 470380 0 180 $X=212840 $Y=464560
X1161 1778 15 14 1026 991 1740 1024 ADDFXL $T=228520 480820 1 180 $X=212840 $Y=480460
X1162 1779 15 14 1060 1064 1739 85 ADDFXL $T=229680 407740 0 180 $X=214000 $Y=401920
X1163 1780 15 14 1071 1015 1770 1029 ADDFXL $T=229680 512140 1 180 $X=214000 $Y=511780
X1164 1781 15 14 615 610 1769 1038 ADDFXL $T=216340 553900 1 0 $X=215740 $Y=548080
X1165 1782 15 14 616 610 1768 1039 ADDFXL $T=216920 543460 1 0 $X=216320 $Y=537640
X1166 1783 15 14 80 1064 1730 99 ADDFXL $T=217500 397300 0 0 $X=216900 $Y=396940
X1167 1784 15 14 1022 951 1697 1042 ADDFXL $T=217500 418180 0 0 $X=216900 $Y=417820
X1168 1785 15 14 612 608 1771 1049 ADDFXL $T=218080 533020 0 0 $X=217480 $Y=532660
X1169 1786 15 14 611 608 1772 1050 ADDFXL $T=218080 543460 0 0 $X=217480 $Y=543100
X1170 1787 15 14 1084 1048 1788 1053 ADDFXL $T=219240 501700 1 0 $X=218640 $Y=495880
X1171 1788 15 14 1072 1015 1773 1028 ADDFXL $T=234320 501700 1 180 $X=218640 $Y=501340
X1172 1789 15 14 1083 1048 1780 1054 ADDFXL $T=219820 512140 1 0 $X=219220 $Y=506320
X1173 1790 15 14 1057 71 1317 101 ADDFXL $T=223880 376420 0 0 $X=223280 $Y=376060
X1174 1791 15 14 1051 963 1778 1065 ADDFXL $T=223880 480820 1 0 $X=223280 $Y=475000
X1175 1792 15 14 1064 979 1776 1058 ADDFXL $T=228520 418180 1 0 $X=227920 $Y=412360
X1176 1793 15 14 1052 963 1777 1066 ADDFXL $T=228520 470380 1 0 $X=227920 $Y=464560
X1177 248 15 14 1094 1080 1779 1055 ADDFXL $T=244760 407740 0 180 $X=229080 $Y=401920
X1178 1794 15 14 1063 979 1784 1059 ADDFXL $T=232580 418180 0 0 $X=231980 $Y=417820
X1179 1795 15 14 1084 1110 1787 1069 ADDFXL $T=249400 501700 0 180 $X=233720 $Y=495880
X1180 1796 15 14 614 612 1782 1074 ADDFXL $T=234320 543460 1 0 $X=233720 $Y=537640
X1181 250 15 14 1095 1080 1783 1056 ADDFXL $T=250560 397300 1 180 $X=234880 $Y=396940
X1182 1159 15 14 613 612 1781 1073 ADDFXL $T=235480 553900 1 0 $X=234880 $Y=548080
X1183 1797 15 14 1110 1019 1775 1078 ADDFXL $T=236060 501700 0 0 $X=235460 $Y=501340
X1184 1168 15 14 1083 1110 1789 1070 ADDFXL $T=251140 512140 0 180 $X=235460 $Y=506320
X1185 1798 15 14 1109 1019 1774 1077 ADDFXL $T=237800 522580 1 0 $X=237200 $Y=516760
X1186 102 15 14 1089 91 1790 107 ADDFXL $T=238960 376420 0 0 $X=238360 $Y=376060
X1187 246 15 14 1067 1007 1791 1081 ADDFXL $T=238960 480820 1 0 $X=238360 $Y=475000
X1188 244 15 14 1068 1007 1793 1082 ADDFXL $T=239540 470380 0 0 $X=238940 $Y=470020
X1189 1799 15 14 1080 983 1792 1090 ADDFXL $T=243600 418180 1 0 $X=243000 $Y=412360
X1190 1762 15 14 1134 1003 1800 1087 ADDFXL $T=244760 407740 1 0 $X=244160 $Y=401920
X1191 1763 15 14 1133 1003 1801 1088 ADDFXL $T=246500 407740 0 0 $X=245900 $Y=407380
X1192 1802 15 14 1079 983 1794 1091 ADDFXL $T=247660 418180 0 0 $X=247060 $Y=417820
X1193 1803 15 14 1120 1037 1797 1104 ADDFXL $T=249400 501700 1 0 $X=248800 $Y=495880
X1194 1804 15 14 618 616 1785 1111 ADDFXL $T=264480 543460 0 180 $X=248800 $Y=537640
X1195 1805 15 14 1119 1037 1798 1103 ADDFXL $T=250560 512140 0 0 $X=249960 $Y=511780
X1196 1800 15 14 1130 987 1799 1117 ADDFXL $T=258680 418180 1 0 $X=258080 $Y=412360
X1197 1801 15 14 1129 987 1802 1118 ADDFXL $T=262740 418180 0 0 $X=262140 $Y=417820
X1198 1806 15 14 1120 1072 1803 1116 ADDFXL $T=264480 501700 1 0 $X=263880 $Y=495880
X1199 1165 15 14 617 616 1786 1112 ADDFXL $T=264480 543460 1 0 $X=263880 $Y=537640
X1200 1163 15 14 1119 1072 1805 1115 ADDFXL $T=265640 512140 0 0 $X=265040 $Y=511780
X1201 562 393 15 14 455 1251 563 1208 1248 OAI222XL $T=465740 522580 1 180 $X=458760 $Y=522220
X1202 1237 15 14 1174 5 234 164 166 161 SDFFRX1 $T=422240 386860 1 0 $X=421640 $Y=381040
X1203 1216 15 14 158 5 165 164 166 169 SDFFRX1 $T=432680 376420 0 0 $X=432080 $Y=376060
X1204 75 80 15 14 1430 78 XOR3XL $T=196040 376420 1 180 $X=178040 $Y=376060
X1205 1106 1068 15 14 1438 1062 XOR3XL $T=250560 459940 0 180 $X=232560 $Y=454120
X1206 1106 1068 15 14 1323 1061 XOR3XL $T=251140 449500 0 180 $X=233140 $Y=443680
X1207 618 614 15 14 1796 1086 XOR3XL $T=235480 533020 0 0 $X=234880 $Y=532660
X1208 1120 1084 15 14 1806 1108 XOR3XL $T=251140 501700 0 0 $X=250540 $Y=501340
X1209 614 618 15 14 1804 1121 XOR3XL $T=256940 533020 0 0 $X=256340 $Y=532660
X1210 1138 1114 15 14 1445 1127 XOR3XL $T=262160 439060 0 0 $X=261560 $Y=438700
X1211 1138 1114 15 14 1331 1128 XOR3XL $T=268540 449500 0 0 $X=267940 $Y=449140
X1212 1084 1120 15 14 1795 1139 XOR3XL $T=268540 501700 0 0 $X=267940 $Y=501340
X1213 1095 1126 15 14 1450 115 XOR3XL $T=305660 386860 0 180 $X=287660 $Y=381040
X1214 1095 1126 15 14 1339 117 XOR3XL $T=310300 376420 1 180 $X=292300 $Y=376060
X1215 739 728 15 14 1252 451 XOR3XL $T=437900 543460 0 0 $X=437300 $Y=543100
X1216 768 728 15 14 1253 460 XOR3XL $T=493000 543460 0 180 $X=475000 $Y=537640
X1217 1611 34 15 14 437 NAND2BX1 $T=50460 386860 1 180 $X=46380 $Y=386500
X1218 1637 469 15 14 492 NAND2BX1 $T=62640 439060 1 180 $X=58560 $Y=438700
X1219 1638 475 15 14 490 NAND2BX1 $T=71920 407740 0 0 $X=71320 $Y=407380
X1220 1652 484 15 14 494 NAND2BX1 $T=89320 459940 0 180 $X=85240 $Y=454120
X1221 1671 499 15 14 509 NAND2BX1 $T=100920 449500 0 180 $X=96840 $Y=443680
X1222 1669 530 15 14 514 NAND2BX1 $T=103240 418180 0 180 $X=99160 $Y=412360
X1223 1666 56 15 14 54 NAND2BX1 $T=116000 386860 1 0 $X=115400 $Y=381040
X1224 1736 540 15 14 538 NAND2BX1 $T=158340 439060 0 180 $X=154260 $Y=433240
X1225 1313 1314 15 14 1551 NAND2BX1 $T=191980 397300 0 180 $X=187900 $Y=391480
X1226 1322 1316 15 14 1554 NAND2BX1 $T=219240 449500 0 0 $X=218640 $Y=449140
X1227 1330 1335 15 14 1557 NAND2BX1 $T=291740 459940 1 180 $X=287660 $Y=459580
X1228 1338 1336 15 14 1560 NAND2BX1 $T=295800 386860 0 0 $X=295200 $Y=386500
X1229 1353 1459 15 14 1491 NAND2BX1 $T=327120 522580 1 180 $X=323040 $Y=522220
X1230 1529 1348 15 14 723 NAND2BX1 $T=332920 480820 1 180 $X=328840 $Y=480460
X1231 1531 1354 15 14 1174 NAND2BX1 $T=346840 418180 0 180 $X=342760 $Y=412360
X1232 330 1293 15 14 1249 NAND2BX1 $T=421080 533020 1 0 $X=420480 $Y=527200
X1233 1293 1304 15 14 798 NAND2BX1 $T=435580 533020 1 0 $X=434980 $Y=527200
X1234 356 1391 15 14 1509 NAND2BX1 $T=446020 522580 1 180 $X=441940 $Y=522220
X1235 1304 1478 15 14 1510 NAND2BX1 $T=446020 522580 0 0 $X=445420 $Y=522220
X1236 1295 1403 15 14 1216 NAND2BX1 $T=481400 428620 1 0 $X=480800 $Y=422800
X1237 1298 1404 15 14 730 NAND2BX1 $T=481980 480820 0 0 $X=481380 $Y=480460
X1238 435 1423 15 14 158 NAND2BX1 $T=528380 407740 1 180 $X=524300 $Y=407380
X1239 797 1264 15 14 1356 556 MX2X1 $T=366560 522580 1 180 $X=360740 $Y=522220
X1240 798 1371 15 14 1266 1198 MX2X1 $T=380480 533020 1 0 $X=379880 $Y=527200
X1241 797 1420 15 14 1418 421 MX2X1 $T=517940 533020 0 180 $X=512120 $Y=527200
X1242 1235 1179 15 14 1236 NAND2XL $T=330600 533020 0 180 $X=327680 $Y=527200
X1243 1262 1232 15 14 1263 NAND2XL $T=531280 533020 1 0 $X=530680 $Y=527200
X1244 1807 15 14 1311 80 1098 AOI2BB1X1 $T=210540 386860 1 180 $X=205300 $Y=386500
X1245 1808 15 14 1320 1068 1105 AOI2BB1X1 $T=244180 459940 1 180 $X=238940 $Y=459580
X1246 1809 15 14 1327 1114 1137 AOI2BB1X1 $T=264480 459940 1 0 $X=263880 $Y=454120
X1247 1810 15 14 1334 1126 1094 AOI2BB1X1 $T=281880 418180 0 180 $X=276640 $Y=412360
X1248 324 15 14 1291 1149 722 AOI2BB1X1 $T=412380 459940 1 180 $X=407140 $Y=459580
X1249 362 15 14 374 737 1216 AOI2BB1X1 $T=440800 418180 1 0 $X=440200 $Y=412360
X1250 358 15 14 368 560 730 AOI2BB1X1 $T=441380 470380 0 0 $X=440780 $Y=470020
X1251 1604 15 14 366 560 731 AOI2BB1X1 $T=447180 480820 1 180 $X=441940 $Y=480460
X1252 1605 15 14 378 737 158 AOI2BB1X1 $T=445440 428620 1 0 $X=444840 $Y=422800
X1253 1811 15 14 1595 792 731 AOI2BB1X1 $T=500540 470380 0 0 $X=499940 $Y=470020
X1254 262 15 14 1238 1237 1349 OAI2BB1X1 $T=341040 407740 1 180 $X=336380 $Y=407380
X1255 272 15 14 1519 646 1237 OAI2BB1X1 $T=354380 397300 0 0 $X=353780 $Y=396940
X1256 374 15 14 1514 158 1395 OAI2BB1X1 $T=454140 418180 1 0 $X=453540 $Y=412360
X1257 1475 15 14 1298 731 1399 OAI2BB1X1 $T=461680 480820 0 0 $X=461080 $Y=480460
X1258 1476 15 14 1295 158 1400 OAI2BB1X1 $T=468640 428620 1 0 $X=468040 $Y=422800
X1259 390 15 14 1517 761 731 OAI2BB1X1 $T=473280 480820 1 0 $X=472680 $Y=475000
X1260 1812 15 14 1421 792 731 OAI2BB1X1 $T=505760 470380 0 180 $X=501100 $Y=464560
X1261 429 15 14 1259 1216 196 OAI2BB1X1 $T=517940 397300 0 0 $X=517340 $Y=396940
X1262 1593 15 14 1261 730 1424 OAI2BB1X1 $T=519680 470380 1 0 $X=519080 $Y=464560
X1263 1579 125 322 15 14 NOR2XL $T=404840 470380 0 0 $X=404240 $Y=470020
X1264 1562 1581 1599 15 14 NOR2XL $T=407160 480820 0 0 $X=406560 $Y=480460
X1265 1582 126 332 15 14 NOR2XL $T=410640 407740 0 0 $X=410040 $Y=407380
X1266 1563 334 1602 15 14 NOR2XL $T=423400 407740 1 180 $X=420480 $Y=407380
X1267 56 15 14 54 1660 AND2X1 $T=113680 386860 0 180 $X=109600 $Y=381040
X1268 62 15 14 56 54 CLKXOR2X1 $T=127600 376420 0 0 $X=127000 $Y=376060
X1269 1807 15 14 1158 1433 1431 NOR3X1 $T=212280 386860 0 0 $X=211680 $Y=386500
X1270 1808 15 14 1161 1440 1439 NOR3X1 $T=245340 459940 0 0 $X=244740 $Y=459580
X1271 1809 15 14 1162 1444 1446 NOR3X1 $T=257520 449500 0 0 $X=256920 $Y=449140
X1272 1810 15 14 1166 1447 1451 NOR3X1 $T=275500 407740 1 180 $X=271420 $Y=407380
X1273 1812 15 14 1526 1811 415 NOR3X1 $T=500540 470380 1 180 $X=496460 $Y=470020
.ends MASCO__P3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cordic_pipeline                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cordic_pipeline GND VDD clk rst theta_in[0] theta_in[10] theta_in[11] theta_in[12] theta_in[13] theta_in[14]
+ theta_in[15] theta_in[1] theta_in[2] theta_in[3] theta_in[4] theta_in[5] theta_in[6] theta_in[7] theta_in[8] theta_in[9]
+ x_in[0] x_in[10] x_in[11] x_in[12] x_in[13] x_in[14] x_in[15] x_in[1] x_in[2] x_in[3]
+ x_in[4] x_in[5] x_in[6] x_in[7] x_in[8] x_in[9] x_out[0] x_out[10] x_out[11] x_out[12]
+ x_out[13] x_out[14] x_out[15] x_out[1] x_out[2] x_out[3] x_out[4] x_out[5] x_out[6] x_out[7]
+ x_out[8] x_out[9] y_in[0] y_in[10] y_in[11] y_in[12] y_in[13] y_in[14] y_in[15] y_in[1]
+ y_in[2] y_in[3] y_in[4] y_in[5] y_in[6] y_in[7] y_in[8] y_in[9] y_out[0] y_out[10]
+ y_out[11] y_out[12] y_out[13] y_out[14] y_out[15] y_out[1] y_out[2] y_out[3] y_out[4] y_out[5]
+ y_out[6] y_out[7] y_out[8] y_out[9]
** N=361 EP=84 FDC=67506
X0 theta_in[13] theta_in[15] theta_in[14] theta_in[7] GND VDD theta_in[8] theta_in[11] theta_in[9] theta_in[12]
+ theta_in[10] theta_in[6] theta_in[4] theta_in[5] clk 23 24 theta_in[3] 26 theta_in[2]
+ 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47
+ 48 49 50 theta_in[1] 52 53 55 56 57 58
+ 59 60 61 62 63 64 65 66 67 68
+ 69 70 71 72 73 74 theta_in[0] 76 77 78
+ 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 96 97 98 99
+ 100 101 102 103 104 106 107 108 109 110
+ 111 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 127 128 129 130 131 132
+ 134 135 136 137 138 140 141 142 143 144
+ 145 146 148 149 150 151 152 153 154 155
+ 156 158 159 160 161 162 163 164 165 167
+ 168 169 170 172 173 174 176 177 178 179
+ 180 181 183 184 185 186 187 188 189 190
+ 191 192 193 194 196 197 198 rst MASCO__P1 $T=0 0 0 0 $X=0 $Y=0
X1 y_in[0] GND VDD x_in[1] 215 216 217 26 218 219
+ clk 30 220 28 221 222 23 24 93 29
+ 72 x_in[2] 62 224 32 38 33 34 35 36
+ 39 37 50 79 42 43 225 226 44 227
+ 64 52 45 47 49 228 229 46 230 48
+ 231 232 53 233 55 59 56 234 235 236
+ 237 60 58 61 238 239 240 41 63 76
+ 65 66 67 77 68 241 69 242 243 244
+ 245 246 73 74 57 247 248 78 249 250
+ 251 252 80 83 81 253 254 84 86 70
+ 90 89 91 88 255 256 257 258 87 259
+ 260 261 262 92 94 263 264 265 266 267
+ 85 268 269 270 271 103 272 273 98 99
+ 71 100 274 101 102 275 276 104 277 106
+ 278 107 110 108 279 280 281 111 282 96
+ 116 97 113 123 114 117 115 125 119 122
+ 124 120 121 137 131 118 127 284 82 285
+ 162 151 286 128 130 129 287 132 148 135
+ 149 138 134 136 109 288 140 143 289 142
+ 290 291 167 141 292 293 144 145 146 152
+ 150 294 153 156 295 296 297 154 298 158
+ 299 155 300 301 159 302 303 165 304 160
+ 161 164 169 170 168 305 192 172 306 173
+ 307 174 308 178 176 309 310 311 179 184
+ 177 187 180 312 185 313 183 314 163 315
+ 316 317 318 319 181 188 320 321 322 323
+ 324 198 191 190 325 326 327 328 329 330
+ 196 331 332 197 MASCO__P2 $T=0 0 0 0 $X=0 $Y=188040
X2 y_in[4] y_in[3] clk y_in[1] y_in[2] GND VDD y_in[11] y_in[7] y_in[8]
+ y_in[6] y_in[5] x_in[3] x_in[5] x_in[6] 23 216 x_in[4] 215 218
+ 222 219 221 x_in[0] 220 x_in[15] x_in[7] 31 224 x_in[8]
+ 40 217 48 x_in[14] 225 241 226 227 64 y_in[9]
+ x_in[9] 229 y_in[12] 228 231 x_in[13] 230 y_in[10] x_in[10] 234
+ 233 237 232 239 238 236 x_in[12] x_in[11] 267 245
+ 243 244 250 246 253 247 248 252 251 249
+ 70 254 263 258 256 255 260 261 275 262
+ 264 259 257 265 242 235 269 y_in[13] 271 272
+ 270 268 273 240 278 276 274 266 277 y_in[15]
+ y_in[14] 279 280 281 282 x_out[13] y_out[4] y_out[8] x_out[15] y_out[6]
+ y_out[5] y_out[7] 189 183 284 y_out[2] 193 y_out[3] 285 y_out[1]
+ 286 y_out[0] 186 287 y_out[9] y_out[10] 290 288 289 x_out[14]
+ x_out[10] y_out[11] y_out[12] y_out[14] x_out[12] y_out[13] 292 296 293 x_out[11]
+ y_out[15] x_out[9] 294 295 297 300 299 309 298 310
+ 301 304 291 303 302 x_out[0] 311 305 307 306
+ x_out[1] x_out[2] 308 316 x_out[8] 312 313 x_out[7] 314 318
+ 317 x_out[6] 321 315 319 x_out[5] 322 324 323 326
+ 320 325 194 330 332 329 327 x_out[3] x_out[4] 328
+ 331 MASCO__P3 $T=0 0 0 0 $X=0 $Y=375960
.ends cordic_pipeline
